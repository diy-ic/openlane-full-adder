magic
tech sky130A
magscale 1 2
timestamp 1702732266
<< viali >>
rect 1409 5661 1443 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 8125 5593 8159 5627
rect 1593 5525 1627 5559
rect 4905 5525 4939 5559
rect 8401 5525 8435 5559
rect 5089 5321 5123 5355
rect 5549 5253 5583 5287
rect 1409 5185 1443 5219
rect 4629 5185 4663 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 8217 5185 8251 5219
rect 4721 5117 4755 5151
rect 5089 5117 5123 5151
rect 4997 5049 5031 5083
rect 1593 4981 1627 5015
rect 5273 4981 5307 5015
rect 8401 4981 8435 5015
rect 4813 4777 4847 4811
rect 4629 4641 4663 4675
rect 1409 4573 1443 4607
rect 4537 4573 4571 4607
rect 1593 4437 1627 4471
<< metal1 >>
rect 1104 7642 8832 7664
rect 1104 7590 2576 7642
rect 2628 7590 2640 7642
rect 2692 7590 2704 7642
rect 2756 7590 2768 7642
rect 2820 7590 2832 7642
rect 2884 7590 4508 7642
rect 4560 7590 4572 7642
rect 4624 7590 4636 7642
rect 4688 7590 4700 7642
rect 4752 7590 4764 7642
rect 4816 7590 6440 7642
rect 6492 7590 6504 7642
rect 6556 7590 6568 7642
rect 6620 7590 6632 7642
rect 6684 7590 6696 7642
rect 6748 7590 8372 7642
rect 8424 7590 8436 7642
rect 8488 7590 8500 7642
rect 8552 7590 8564 7642
rect 8616 7590 8628 7642
rect 8680 7590 8832 7642
rect 1104 7568 8832 7590
rect 1104 7098 8832 7120
rect 1104 7046 1916 7098
rect 1968 7046 1980 7098
rect 2032 7046 2044 7098
rect 2096 7046 2108 7098
rect 2160 7046 2172 7098
rect 2224 7046 3848 7098
rect 3900 7046 3912 7098
rect 3964 7046 3976 7098
rect 4028 7046 4040 7098
rect 4092 7046 4104 7098
rect 4156 7046 5780 7098
rect 5832 7046 5844 7098
rect 5896 7046 5908 7098
rect 5960 7046 5972 7098
rect 6024 7046 6036 7098
rect 6088 7046 7712 7098
rect 7764 7046 7776 7098
rect 7828 7046 7840 7098
rect 7892 7046 7904 7098
rect 7956 7046 7968 7098
rect 8020 7046 8832 7098
rect 1104 7024 8832 7046
rect 1104 6554 8832 6576
rect 1104 6502 2576 6554
rect 2628 6502 2640 6554
rect 2692 6502 2704 6554
rect 2756 6502 2768 6554
rect 2820 6502 2832 6554
rect 2884 6502 4508 6554
rect 4560 6502 4572 6554
rect 4624 6502 4636 6554
rect 4688 6502 4700 6554
rect 4752 6502 4764 6554
rect 4816 6502 6440 6554
rect 6492 6502 6504 6554
rect 6556 6502 6568 6554
rect 6620 6502 6632 6554
rect 6684 6502 6696 6554
rect 6748 6502 8372 6554
rect 8424 6502 8436 6554
rect 8488 6502 8500 6554
rect 8552 6502 8564 6554
rect 8616 6502 8628 6554
rect 8680 6502 8832 6554
rect 1104 6480 8832 6502
rect 1104 6010 8832 6032
rect 1104 5958 1916 6010
rect 1968 5958 1980 6010
rect 2032 5958 2044 6010
rect 2096 5958 2108 6010
rect 2160 5958 2172 6010
rect 2224 5958 3848 6010
rect 3900 5958 3912 6010
rect 3964 5958 3976 6010
rect 4028 5958 4040 6010
rect 4092 5958 4104 6010
rect 4156 5958 5780 6010
rect 5832 5958 5844 6010
rect 5896 5958 5908 6010
rect 5960 5958 5972 6010
rect 6024 5958 6036 6010
rect 6088 5958 7712 6010
rect 7764 5958 7776 6010
rect 7828 5958 7840 6010
rect 7892 5958 7904 6010
rect 7956 5958 7968 6010
rect 8020 5958 8832 6010
rect 1104 5936 8832 5958
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4304 5732 4936 5760
rect 4304 5720 4310 5732
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 4908 5701 4936 5732
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4448 5664 4721 5692
rect 4448 5568 4476 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 8110 5584 8116 5636
rect 8168 5584 8174 5636
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 4154 5556 4160 5568
rect 1627 5528 4160 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4430 5516 4436 5568
rect 4488 5516 4494 5568
rect 4890 5516 4896 5568
rect 4948 5516 4954 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 8754 5556 8760 5568
rect 8435 5528 8760 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 1104 5466 8832 5488
rect 1104 5414 2576 5466
rect 2628 5414 2640 5466
rect 2692 5414 2704 5466
rect 2756 5414 2768 5466
rect 2820 5414 2832 5466
rect 2884 5414 4508 5466
rect 4560 5414 4572 5466
rect 4624 5414 4636 5466
rect 4688 5414 4700 5466
rect 4752 5414 4764 5466
rect 4816 5414 6440 5466
rect 6492 5414 6504 5466
rect 6556 5414 6568 5466
rect 6620 5414 6632 5466
rect 6684 5414 6696 5466
rect 6748 5414 8372 5466
rect 8424 5414 8436 5466
rect 8488 5414 8500 5466
rect 8552 5414 8564 5466
rect 8616 5414 8628 5466
rect 8680 5414 8832 5466
rect 1104 5392 8832 5414
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 8110 5352 8116 5364
rect 5123 5324 8116 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 5368 5256 5549 5284
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 5368 5225 5396 5256
rect 5537 5253 5549 5256
rect 5583 5253 5595 5287
rect 5537 5247 5595 5253
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4212 5188 4629 5216
rect 4212 5176 4218 5188
rect 4617 5185 4629 5188
rect 4663 5216 4675 5219
rect 5353 5219 5411 5225
rect 4663 5188 5304 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4755 5120 4844 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 4246 5012 4252 5024
rect 1627 4984 4252 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4816 5012 4844 5120
rect 4890 5108 4896 5160
rect 4948 5148 4954 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4948 5120 5089 5148
rect 4948 5108 4954 5120
rect 5077 5117 5089 5120
rect 5123 5117 5135 5151
rect 5276 5148 5304 5188
rect 5353 5185 5365 5219
rect 5399 5185 5411 5219
rect 5353 5179 5411 5185
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 5445 5179 5503 5185
rect 6886 5188 8217 5216
rect 5460 5148 5488 5179
rect 5276 5120 5488 5148
rect 5077 5111 5135 5117
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 6886 5080 6914 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 5031 5052 6914 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 4890 5012 4896 5024
rect 4816 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 5012 4954 5024
rect 5261 5015 5319 5021
rect 5261 5012 5273 5015
rect 4948 4984 5273 5012
rect 4948 4972 4954 4984
rect 5261 4981 5273 4984
rect 5307 4981 5319 5015
rect 5261 4975 5319 4981
rect 8386 4972 8392 5024
rect 8444 4972 8450 5024
rect 1104 4922 8832 4944
rect 1104 4870 1916 4922
rect 1968 4870 1980 4922
rect 2032 4870 2044 4922
rect 2096 4870 2108 4922
rect 2160 4870 2172 4922
rect 2224 4870 3848 4922
rect 3900 4870 3912 4922
rect 3964 4870 3976 4922
rect 4028 4870 4040 4922
rect 4092 4870 4104 4922
rect 4156 4870 5780 4922
rect 5832 4870 5844 4922
rect 5896 4870 5908 4922
rect 5960 4870 5972 4922
rect 6024 4870 6036 4922
rect 6088 4870 7712 4922
rect 7764 4870 7776 4922
rect 7828 4870 7840 4922
rect 7892 4870 7904 4922
rect 7956 4870 7968 4922
rect 8020 4870 8832 4922
rect 1104 4848 8832 4870
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4808 4859 4811
rect 4890 4808 4896 4820
rect 4847 4780 4896 4808
rect 4847 4777 4859 4780
rect 4801 4771 4859 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 4246 4564 4252 4616
rect 4304 4604 4310 4616
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 4304 4576 4537 4604
rect 4304 4564 4310 4576
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 4430 4468 4436 4480
rect 1627 4440 4436 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 4430 4428 4436 4440
rect 4488 4468 4494 4480
rect 4632 4468 4660 4635
rect 4488 4440 4660 4468
rect 4488 4428 4494 4440
rect 1104 4378 8832 4400
rect 1104 4326 2576 4378
rect 2628 4326 2640 4378
rect 2692 4326 2704 4378
rect 2756 4326 2768 4378
rect 2820 4326 2832 4378
rect 2884 4326 4508 4378
rect 4560 4326 4572 4378
rect 4624 4326 4636 4378
rect 4688 4326 4700 4378
rect 4752 4326 4764 4378
rect 4816 4326 6440 4378
rect 6492 4326 6504 4378
rect 6556 4326 6568 4378
rect 6620 4326 6632 4378
rect 6684 4326 6696 4378
rect 6748 4326 8372 4378
rect 8424 4326 8436 4378
rect 8488 4326 8500 4378
rect 8552 4326 8564 4378
rect 8616 4326 8628 4378
rect 8680 4326 8832 4378
rect 1104 4304 8832 4326
rect 1104 3834 8832 3856
rect 1104 3782 1916 3834
rect 1968 3782 1980 3834
rect 2032 3782 2044 3834
rect 2096 3782 2108 3834
rect 2160 3782 2172 3834
rect 2224 3782 3848 3834
rect 3900 3782 3912 3834
rect 3964 3782 3976 3834
rect 4028 3782 4040 3834
rect 4092 3782 4104 3834
rect 4156 3782 5780 3834
rect 5832 3782 5844 3834
rect 5896 3782 5908 3834
rect 5960 3782 5972 3834
rect 6024 3782 6036 3834
rect 6088 3782 7712 3834
rect 7764 3782 7776 3834
rect 7828 3782 7840 3834
rect 7892 3782 7904 3834
rect 7956 3782 7968 3834
rect 8020 3782 8832 3834
rect 1104 3760 8832 3782
rect 1104 3290 8832 3312
rect 1104 3238 2576 3290
rect 2628 3238 2640 3290
rect 2692 3238 2704 3290
rect 2756 3238 2768 3290
rect 2820 3238 2832 3290
rect 2884 3238 4508 3290
rect 4560 3238 4572 3290
rect 4624 3238 4636 3290
rect 4688 3238 4700 3290
rect 4752 3238 4764 3290
rect 4816 3238 6440 3290
rect 6492 3238 6504 3290
rect 6556 3238 6568 3290
rect 6620 3238 6632 3290
rect 6684 3238 6696 3290
rect 6748 3238 8372 3290
rect 8424 3238 8436 3290
rect 8488 3238 8500 3290
rect 8552 3238 8564 3290
rect 8616 3238 8628 3290
rect 8680 3238 8832 3290
rect 1104 3216 8832 3238
rect 1104 2746 8832 2768
rect 1104 2694 1916 2746
rect 1968 2694 1980 2746
rect 2032 2694 2044 2746
rect 2096 2694 2108 2746
rect 2160 2694 2172 2746
rect 2224 2694 3848 2746
rect 3900 2694 3912 2746
rect 3964 2694 3976 2746
rect 4028 2694 4040 2746
rect 4092 2694 4104 2746
rect 4156 2694 5780 2746
rect 5832 2694 5844 2746
rect 5896 2694 5908 2746
rect 5960 2694 5972 2746
rect 6024 2694 6036 2746
rect 6088 2694 7712 2746
rect 7764 2694 7776 2746
rect 7828 2694 7840 2746
rect 7892 2694 7904 2746
rect 7956 2694 7968 2746
rect 8020 2694 8832 2746
rect 1104 2672 8832 2694
rect 1104 2202 8832 2224
rect 1104 2150 2576 2202
rect 2628 2150 2640 2202
rect 2692 2150 2704 2202
rect 2756 2150 2768 2202
rect 2820 2150 2832 2202
rect 2884 2150 4508 2202
rect 4560 2150 4572 2202
rect 4624 2150 4636 2202
rect 4688 2150 4700 2202
rect 4752 2150 4764 2202
rect 4816 2150 6440 2202
rect 6492 2150 6504 2202
rect 6556 2150 6568 2202
rect 6620 2150 6632 2202
rect 6684 2150 6696 2202
rect 6748 2150 8372 2202
rect 8424 2150 8436 2202
rect 8488 2150 8500 2202
rect 8552 2150 8564 2202
rect 8616 2150 8628 2202
rect 8680 2150 8832 2202
rect 1104 2128 8832 2150
<< via1 >>
rect 2576 7590 2628 7642
rect 2640 7590 2692 7642
rect 2704 7590 2756 7642
rect 2768 7590 2820 7642
rect 2832 7590 2884 7642
rect 4508 7590 4560 7642
rect 4572 7590 4624 7642
rect 4636 7590 4688 7642
rect 4700 7590 4752 7642
rect 4764 7590 4816 7642
rect 6440 7590 6492 7642
rect 6504 7590 6556 7642
rect 6568 7590 6620 7642
rect 6632 7590 6684 7642
rect 6696 7590 6748 7642
rect 8372 7590 8424 7642
rect 8436 7590 8488 7642
rect 8500 7590 8552 7642
rect 8564 7590 8616 7642
rect 8628 7590 8680 7642
rect 1916 7046 1968 7098
rect 1980 7046 2032 7098
rect 2044 7046 2096 7098
rect 2108 7046 2160 7098
rect 2172 7046 2224 7098
rect 3848 7046 3900 7098
rect 3912 7046 3964 7098
rect 3976 7046 4028 7098
rect 4040 7046 4092 7098
rect 4104 7046 4156 7098
rect 5780 7046 5832 7098
rect 5844 7046 5896 7098
rect 5908 7046 5960 7098
rect 5972 7046 6024 7098
rect 6036 7046 6088 7098
rect 7712 7046 7764 7098
rect 7776 7046 7828 7098
rect 7840 7046 7892 7098
rect 7904 7046 7956 7098
rect 7968 7046 8020 7098
rect 2576 6502 2628 6554
rect 2640 6502 2692 6554
rect 2704 6502 2756 6554
rect 2768 6502 2820 6554
rect 2832 6502 2884 6554
rect 4508 6502 4560 6554
rect 4572 6502 4624 6554
rect 4636 6502 4688 6554
rect 4700 6502 4752 6554
rect 4764 6502 4816 6554
rect 6440 6502 6492 6554
rect 6504 6502 6556 6554
rect 6568 6502 6620 6554
rect 6632 6502 6684 6554
rect 6696 6502 6748 6554
rect 8372 6502 8424 6554
rect 8436 6502 8488 6554
rect 8500 6502 8552 6554
rect 8564 6502 8616 6554
rect 8628 6502 8680 6554
rect 1916 5958 1968 6010
rect 1980 5958 2032 6010
rect 2044 5958 2096 6010
rect 2108 5958 2160 6010
rect 2172 5958 2224 6010
rect 3848 5958 3900 6010
rect 3912 5958 3964 6010
rect 3976 5958 4028 6010
rect 4040 5958 4092 6010
rect 4104 5958 4156 6010
rect 5780 5958 5832 6010
rect 5844 5958 5896 6010
rect 5908 5958 5960 6010
rect 5972 5958 6024 6010
rect 6036 5958 6088 6010
rect 7712 5958 7764 6010
rect 7776 5958 7828 6010
rect 7840 5958 7892 6010
rect 7904 5958 7956 6010
rect 7968 5958 8020 6010
rect 4252 5720 4304 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 8116 5627 8168 5636
rect 8116 5593 8125 5627
rect 8125 5593 8159 5627
rect 8159 5593 8168 5627
rect 8116 5584 8168 5593
rect 4160 5516 4212 5568
rect 4436 5516 4488 5568
rect 4896 5559 4948 5568
rect 4896 5525 4905 5559
rect 4905 5525 4939 5559
rect 4939 5525 4948 5559
rect 4896 5516 4948 5525
rect 8760 5516 8812 5568
rect 2576 5414 2628 5466
rect 2640 5414 2692 5466
rect 2704 5414 2756 5466
rect 2768 5414 2820 5466
rect 2832 5414 2884 5466
rect 4508 5414 4560 5466
rect 4572 5414 4624 5466
rect 4636 5414 4688 5466
rect 4700 5414 4752 5466
rect 4764 5414 4816 5466
rect 6440 5414 6492 5466
rect 6504 5414 6556 5466
rect 6568 5414 6620 5466
rect 6632 5414 6684 5466
rect 6696 5414 6748 5466
rect 8372 5414 8424 5466
rect 8436 5414 8488 5466
rect 8500 5414 8552 5466
rect 8564 5414 8616 5466
rect 8628 5414 8680 5466
rect 8116 5312 8168 5364
rect 940 5176 992 5228
rect 4160 5176 4212 5228
rect 4252 4972 4304 5024
rect 4896 5108 4948 5160
rect 4896 4972 4948 5024
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 1916 4870 1968 4922
rect 1980 4870 2032 4922
rect 2044 4870 2096 4922
rect 2108 4870 2160 4922
rect 2172 4870 2224 4922
rect 3848 4870 3900 4922
rect 3912 4870 3964 4922
rect 3976 4870 4028 4922
rect 4040 4870 4092 4922
rect 4104 4870 4156 4922
rect 5780 4870 5832 4922
rect 5844 4870 5896 4922
rect 5908 4870 5960 4922
rect 5972 4870 6024 4922
rect 6036 4870 6088 4922
rect 7712 4870 7764 4922
rect 7776 4870 7828 4922
rect 7840 4870 7892 4922
rect 7904 4870 7956 4922
rect 7968 4870 8020 4922
rect 4896 4768 4948 4820
rect 940 4564 992 4616
rect 4252 4564 4304 4616
rect 4436 4428 4488 4480
rect 2576 4326 2628 4378
rect 2640 4326 2692 4378
rect 2704 4326 2756 4378
rect 2768 4326 2820 4378
rect 2832 4326 2884 4378
rect 4508 4326 4560 4378
rect 4572 4326 4624 4378
rect 4636 4326 4688 4378
rect 4700 4326 4752 4378
rect 4764 4326 4816 4378
rect 6440 4326 6492 4378
rect 6504 4326 6556 4378
rect 6568 4326 6620 4378
rect 6632 4326 6684 4378
rect 6696 4326 6748 4378
rect 8372 4326 8424 4378
rect 8436 4326 8488 4378
rect 8500 4326 8552 4378
rect 8564 4326 8616 4378
rect 8628 4326 8680 4378
rect 1916 3782 1968 3834
rect 1980 3782 2032 3834
rect 2044 3782 2096 3834
rect 2108 3782 2160 3834
rect 2172 3782 2224 3834
rect 3848 3782 3900 3834
rect 3912 3782 3964 3834
rect 3976 3782 4028 3834
rect 4040 3782 4092 3834
rect 4104 3782 4156 3834
rect 5780 3782 5832 3834
rect 5844 3782 5896 3834
rect 5908 3782 5960 3834
rect 5972 3782 6024 3834
rect 6036 3782 6088 3834
rect 7712 3782 7764 3834
rect 7776 3782 7828 3834
rect 7840 3782 7892 3834
rect 7904 3782 7956 3834
rect 7968 3782 8020 3834
rect 2576 3238 2628 3290
rect 2640 3238 2692 3290
rect 2704 3238 2756 3290
rect 2768 3238 2820 3290
rect 2832 3238 2884 3290
rect 4508 3238 4560 3290
rect 4572 3238 4624 3290
rect 4636 3238 4688 3290
rect 4700 3238 4752 3290
rect 4764 3238 4816 3290
rect 6440 3238 6492 3290
rect 6504 3238 6556 3290
rect 6568 3238 6620 3290
rect 6632 3238 6684 3290
rect 6696 3238 6748 3290
rect 8372 3238 8424 3290
rect 8436 3238 8488 3290
rect 8500 3238 8552 3290
rect 8564 3238 8616 3290
rect 8628 3238 8680 3290
rect 1916 2694 1968 2746
rect 1980 2694 2032 2746
rect 2044 2694 2096 2746
rect 2108 2694 2160 2746
rect 2172 2694 2224 2746
rect 3848 2694 3900 2746
rect 3912 2694 3964 2746
rect 3976 2694 4028 2746
rect 4040 2694 4092 2746
rect 4104 2694 4156 2746
rect 5780 2694 5832 2746
rect 5844 2694 5896 2746
rect 5908 2694 5960 2746
rect 5972 2694 6024 2746
rect 6036 2694 6088 2746
rect 7712 2694 7764 2746
rect 7776 2694 7828 2746
rect 7840 2694 7892 2746
rect 7904 2694 7956 2746
rect 7968 2694 8020 2746
rect 2576 2150 2628 2202
rect 2640 2150 2692 2202
rect 2704 2150 2756 2202
rect 2768 2150 2820 2202
rect 2832 2150 2884 2202
rect 4508 2150 4560 2202
rect 4572 2150 4624 2202
rect 4636 2150 4688 2202
rect 4700 2150 4752 2202
rect 4764 2150 4816 2202
rect 6440 2150 6492 2202
rect 6504 2150 6556 2202
rect 6568 2150 6620 2202
rect 6632 2150 6684 2202
rect 6696 2150 6748 2202
rect 8372 2150 8424 2202
rect 8436 2150 8488 2202
rect 8500 2150 8552 2202
rect 8564 2150 8616 2202
rect 8628 2150 8680 2202
<< metal2 >>
rect 2576 7644 2884 7653
rect 2576 7642 2582 7644
rect 2638 7642 2662 7644
rect 2718 7642 2742 7644
rect 2798 7642 2822 7644
rect 2878 7642 2884 7644
rect 2638 7590 2640 7642
rect 2820 7590 2822 7642
rect 2576 7588 2582 7590
rect 2638 7588 2662 7590
rect 2718 7588 2742 7590
rect 2798 7588 2822 7590
rect 2878 7588 2884 7590
rect 2576 7579 2884 7588
rect 4508 7644 4816 7653
rect 4508 7642 4514 7644
rect 4570 7642 4594 7644
rect 4650 7642 4674 7644
rect 4730 7642 4754 7644
rect 4810 7642 4816 7644
rect 4570 7590 4572 7642
rect 4752 7590 4754 7642
rect 4508 7588 4514 7590
rect 4570 7588 4594 7590
rect 4650 7588 4674 7590
rect 4730 7588 4754 7590
rect 4810 7588 4816 7590
rect 4508 7579 4816 7588
rect 6440 7644 6748 7653
rect 6440 7642 6446 7644
rect 6502 7642 6526 7644
rect 6582 7642 6606 7644
rect 6662 7642 6686 7644
rect 6742 7642 6748 7644
rect 6502 7590 6504 7642
rect 6684 7590 6686 7642
rect 6440 7588 6446 7590
rect 6502 7588 6526 7590
rect 6582 7588 6606 7590
rect 6662 7588 6686 7590
rect 6742 7588 6748 7590
rect 6440 7579 6748 7588
rect 8372 7644 8680 7653
rect 8372 7642 8378 7644
rect 8434 7642 8458 7644
rect 8514 7642 8538 7644
rect 8594 7642 8618 7644
rect 8674 7642 8680 7644
rect 8434 7590 8436 7642
rect 8616 7590 8618 7642
rect 8372 7588 8378 7590
rect 8434 7588 8458 7590
rect 8514 7588 8538 7590
rect 8594 7588 8618 7590
rect 8674 7588 8680 7590
rect 8372 7579 8680 7588
rect 1916 7100 2224 7109
rect 1916 7098 1922 7100
rect 1978 7098 2002 7100
rect 2058 7098 2082 7100
rect 2138 7098 2162 7100
rect 2218 7098 2224 7100
rect 1978 7046 1980 7098
rect 2160 7046 2162 7098
rect 1916 7044 1922 7046
rect 1978 7044 2002 7046
rect 2058 7044 2082 7046
rect 2138 7044 2162 7046
rect 2218 7044 2224 7046
rect 1916 7035 2224 7044
rect 3848 7100 4156 7109
rect 3848 7098 3854 7100
rect 3910 7098 3934 7100
rect 3990 7098 4014 7100
rect 4070 7098 4094 7100
rect 4150 7098 4156 7100
rect 3910 7046 3912 7098
rect 4092 7046 4094 7098
rect 3848 7044 3854 7046
rect 3910 7044 3934 7046
rect 3990 7044 4014 7046
rect 4070 7044 4094 7046
rect 4150 7044 4156 7046
rect 3848 7035 4156 7044
rect 5780 7100 6088 7109
rect 5780 7098 5786 7100
rect 5842 7098 5866 7100
rect 5922 7098 5946 7100
rect 6002 7098 6026 7100
rect 6082 7098 6088 7100
rect 5842 7046 5844 7098
rect 6024 7046 6026 7098
rect 5780 7044 5786 7046
rect 5842 7044 5866 7046
rect 5922 7044 5946 7046
rect 6002 7044 6026 7046
rect 6082 7044 6088 7046
rect 5780 7035 6088 7044
rect 7712 7100 8020 7109
rect 7712 7098 7718 7100
rect 7774 7098 7798 7100
rect 7854 7098 7878 7100
rect 7934 7098 7958 7100
rect 8014 7098 8020 7100
rect 7774 7046 7776 7098
rect 7956 7046 7958 7098
rect 7712 7044 7718 7046
rect 7774 7044 7798 7046
rect 7854 7044 7878 7046
rect 7934 7044 7958 7046
rect 8014 7044 8020 7046
rect 7712 7035 8020 7044
rect 2576 6556 2884 6565
rect 2576 6554 2582 6556
rect 2638 6554 2662 6556
rect 2718 6554 2742 6556
rect 2798 6554 2822 6556
rect 2878 6554 2884 6556
rect 2638 6502 2640 6554
rect 2820 6502 2822 6554
rect 2576 6500 2582 6502
rect 2638 6500 2662 6502
rect 2718 6500 2742 6502
rect 2798 6500 2822 6502
rect 2878 6500 2884 6502
rect 2576 6491 2884 6500
rect 4508 6556 4816 6565
rect 4508 6554 4514 6556
rect 4570 6554 4594 6556
rect 4650 6554 4674 6556
rect 4730 6554 4754 6556
rect 4810 6554 4816 6556
rect 4570 6502 4572 6554
rect 4752 6502 4754 6554
rect 4508 6500 4514 6502
rect 4570 6500 4594 6502
rect 4650 6500 4674 6502
rect 4730 6500 4754 6502
rect 4810 6500 4816 6502
rect 4508 6491 4816 6500
rect 6440 6556 6748 6565
rect 6440 6554 6446 6556
rect 6502 6554 6526 6556
rect 6582 6554 6606 6556
rect 6662 6554 6686 6556
rect 6742 6554 6748 6556
rect 6502 6502 6504 6554
rect 6684 6502 6686 6554
rect 6440 6500 6446 6502
rect 6502 6500 6526 6502
rect 6582 6500 6606 6502
rect 6662 6500 6686 6502
rect 6742 6500 6748 6502
rect 6440 6491 6748 6500
rect 8372 6556 8680 6565
rect 8372 6554 8378 6556
rect 8434 6554 8458 6556
rect 8514 6554 8538 6556
rect 8594 6554 8618 6556
rect 8674 6554 8680 6556
rect 8434 6502 8436 6554
rect 8616 6502 8618 6554
rect 8372 6500 8378 6502
rect 8434 6500 8458 6502
rect 8514 6500 8538 6502
rect 8594 6500 8618 6502
rect 8674 6500 8680 6502
rect 8372 6491 8680 6500
rect 1916 6012 2224 6021
rect 1916 6010 1922 6012
rect 1978 6010 2002 6012
rect 2058 6010 2082 6012
rect 2138 6010 2162 6012
rect 2218 6010 2224 6012
rect 1978 5958 1980 6010
rect 2160 5958 2162 6010
rect 1916 5956 1922 5958
rect 1978 5956 2002 5958
rect 2058 5956 2082 5958
rect 2138 5956 2162 5958
rect 2218 5956 2224 5958
rect 1916 5947 2224 5956
rect 3848 6012 4156 6021
rect 3848 6010 3854 6012
rect 3910 6010 3934 6012
rect 3990 6010 4014 6012
rect 4070 6010 4094 6012
rect 4150 6010 4156 6012
rect 3910 5958 3912 6010
rect 4092 5958 4094 6010
rect 3848 5956 3854 5958
rect 3910 5956 3934 5958
rect 3990 5956 4014 5958
rect 4070 5956 4094 5958
rect 4150 5956 4156 5958
rect 3848 5947 4156 5956
rect 5780 6012 6088 6021
rect 5780 6010 5786 6012
rect 5842 6010 5866 6012
rect 5922 6010 5946 6012
rect 6002 6010 6026 6012
rect 6082 6010 6088 6012
rect 5842 5958 5844 6010
rect 6024 5958 6026 6010
rect 5780 5956 5786 5958
rect 5842 5956 5866 5958
rect 5922 5956 5946 5958
rect 6002 5956 6026 5958
rect 6082 5956 6088 5958
rect 5780 5947 6088 5956
rect 7712 6012 8020 6021
rect 7712 6010 7718 6012
rect 7774 6010 7798 6012
rect 7854 6010 7878 6012
rect 7934 6010 7958 6012
rect 8014 6010 8020 6012
rect 7774 5958 7776 6010
rect 7956 5958 7958 6010
rect 7712 5956 7718 5958
rect 7774 5956 7798 5958
rect 7854 5956 7878 5958
rect 7934 5956 7958 5958
rect 8014 5956 8020 5958
rect 7712 5947 8020 5956
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 4160 5568 4212 5574
rect 1398 5536 1454 5545
rect 4160 5510 4212 5516
rect 1398 5471 1454 5480
rect 2576 5468 2884 5477
rect 2576 5466 2582 5468
rect 2638 5466 2662 5468
rect 2718 5466 2742 5468
rect 2798 5466 2822 5468
rect 2878 5466 2884 5468
rect 2638 5414 2640 5466
rect 2820 5414 2822 5466
rect 2576 5412 2582 5414
rect 2638 5412 2662 5414
rect 2718 5412 2742 5414
rect 2798 5412 2822 5414
rect 2878 5412 2884 5414
rect 2576 5403 2884 5412
rect 4172 5234 4200 5510
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 952 4865 980 5170
rect 4264 5030 4292 5714
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 1916 4924 2224 4933
rect 1916 4922 1922 4924
rect 1978 4922 2002 4924
rect 2058 4922 2082 4924
rect 2138 4922 2162 4924
rect 2218 4922 2224 4924
rect 1978 4870 1980 4922
rect 2160 4870 2162 4922
rect 1916 4868 1922 4870
rect 1978 4868 2002 4870
rect 2058 4868 2082 4870
rect 2138 4868 2162 4870
rect 2218 4868 2224 4870
rect 938 4856 994 4865
rect 1916 4859 2224 4868
rect 3848 4924 4156 4933
rect 3848 4922 3854 4924
rect 3910 4922 3934 4924
rect 3990 4922 4014 4924
rect 4070 4922 4094 4924
rect 4150 4922 4156 4924
rect 3910 4870 3912 4922
rect 4092 4870 4094 4922
rect 3848 4868 3854 4870
rect 3910 4868 3934 4870
rect 3990 4868 4014 4870
rect 4070 4868 4094 4870
rect 4150 4868 4156 4870
rect 3848 4859 4156 4868
rect 938 4791 994 4800
rect 4264 4622 4292 4966
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 952 4185 980 4558
rect 4448 4486 4476 5510
rect 4508 5468 4816 5477
rect 4508 5466 4514 5468
rect 4570 5466 4594 5468
rect 4650 5466 4674 5468
rect 4730 5466 4754 5468
rect 4810 5466 4816 5468
rect 4570 5414 4572 5466
rect 4752 5414 4754 5466
rect 4508 5412 4514 5414
rect 4570 5412 4594 5414
rect 4650 5412 4674 5414
rect 4730 5412 4754 5414
rect 4810 5412 4816 5414
rect 4508 5403 4816 5412
rect 4908 5166 4936 5510
rect 6440 5468 6748 5477
rect 6440 5466 6446 5468
rect 6502 5466 6526 5468
rect 6582 5466 6606 5468
rect 6662 5466 6686 5468
rect 6742 5466 6748 5468
rect 6502 5414 6504 5466
rect 6684 5414 6686 5466
rect 6440 5412 6446 5414
rect 6502 5412 6526 5414
rect 6582 5412 6606 5414
rect 6662 5412 6686 5414
rect 6742 5412 6748 5414
rect 6440 5403 6748 5412
rect 8128 5370 8156 5578
rect 8760 5568 8812 5574
rect 8758 5536 8760 5545
rect 8812 5536 8814 5545
rect 8372 5468 8680 5477
rect 8758 5471 8814 5480
rect 8372 5466 8378 5468
rect 8434 5466 8458 5468
rect 8514 5466 8538 5468
rect 8594 5466 8618 5468
rect 8674 5466 8680 5468
rect 8434 5414 8436 5466
rect 8616 5414 8618 5466
rect 8372 5412 8378 5414
rect 8434 5412 8458 5414
rect 8514 5412 8538 5414
rect 8594 5412 8618 5414
rect 8674 5412 8680 5414
rect 8372 5403 8680 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 4908 4826 4936 4966
rect 5780 4924 6088 4933
rect 5780 4922 5786 4924
rect 5842 4922 5866 4924
rect 5922 4922 5946 4924
rect 6002 4922 6026 4924
rect 6082 4922 6088 4924
rect 5842 4870 5844 4922
rect 6024 4870 6026 4922
rect 5780 4868 5786 4870
rect 5842 4868 5866 4870
rect 5922 4868 5946 4870
rect 6002 4868 6026 4870
rect 6082 4868 6088 4870
rect 5780 4859 6088 4868
rect 7712 4924 8020 4933
rect 7712 4922 7718 4924
rect 7774 4922 7798 4924
rect 7854 4922 7878 4924
rect 7934 4922 7958 4924
rect 8014 4922 8020 4924
rect 7774 4870 7776 4922
rect 7956 4870 7958 4922
rect 7712 4868 7718 4870
rect 7774 4868 7798 4870
rect 7854 4868 7878 4870
rect 7934 4868 7958 4870
rect 8014 4868 8020 4870
rect 7712 4859 8020 4868
rect 8404 4865 8432 4966
rect 8390 4856 8446 4865
rect 4896 4820 4948 4826
rect 8390 4791 8446 4800
rect 4896 4762 4948 4768
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 2576 4380 2884 4389
rect 2576 4378 2582 4380
rect 2638 4378 2662 4380
rect 2718 4378 2742 4380
rect 2798 4378 2822 4380
rect 2878 4378 2884 4380
rect 2638 4326 2640 4378
rect 2820 4326 2822 4378
rect 2576 4324 2582 4326
rect 2638 4324 2662 4326
rect 2718 4324 2742 4326
rect 2798 4324 2822 4326
rect 2878 4324 2884 4326
rect 2576 4315 2884 4324
rect 4508 4380 4816 4389
rect 4508 4378 4514 4380
rect 4570 4378 4594 4380
rect 4650 4378 4674 4380
rect 4730 4378 4754 4380
rect 4810 4378 4816 4380
rect 4570 4326 4572 4378
rect 4752 4326 4754 4378
rect 4508 4324 4514 4326
rect 4570 4324 4594 4326
rect 4650 4324 4674 4326
rect 4730 4324 4754 4326
rect 4810 4324 4816 4326
rect 4508 4315 4816 4324
rect 6440 4380 6748 4389
rect 6440 4378 6446 4380
rect 6502 4378 6526 4380
rect 6582 4378 6606 4380
rect 6662 4378 6686 4380
rect 6742 4378 6748 4380
rect 6502 4326 6504 4378
rect 6684 4326 6686 4378
rect 6440 4324 6446 4326
rect 6502 4324 6526 4326
rect 6582 4324 6606 4326
rect 6662 4324 6686 4326
rect 6742 4324 6748 4326
rect 6440 4315 6748 4324
rect 8372 4380 8680 4389
rect 8372 4378 8378 4380
rect 8434 4378 8458 4380
rect 8514 4378 8538 4380
rect 8594 4378 8618 4380
rect 8674 4378 8680 4380
rect 8434 4326 8436 4378
rect 8616 4326 8618 4378
rect 8372 4324 8378 4326
rect 8434 4324 8458 4326
rect 8514 4324 8538 4326
rect 8594 4324 8618 4326
rect 8674 4324 8680 4326
rect 8372 4315 8680 4324
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1916 3836 2224 3845
rect 1916 3834 1922 3836
rect 1978 3834 2002 3836
rect 2058 3834 2082 3836
rect 2138 3834 2162 3836
rect 2218 3834 2224 3836
rect 1978 3782 1980 3834
rect 2160 3782 2162 3834
rect 1916 3780 1922 3782
rect 1978 3780 2002 3782
rect 2058 3780 2082 3782
rect 2138 3780 2162 3782
rect 2218 3780 2224 3782
rect 1916 3771 2224 3780
rect 3848 3836 4156 3845
rect 3848 3834 3854 3836
rect 3910 3834 3934 3836
rect 3990 3834 4014 3836
rect 4070 3834 4094 3836
rect 4150 3834 4156 3836
rect 3910 3782 3912 3834
rect 4092 3782 4094 3834
rect 3848 3780 3854 3782
rect 3910 3780 3934 3782
rect 3990 3780 4014 3782
rect 4070 3780 4094 3782
rect 4150 3780 4156 3782
rect 3848 3771 4156 3780
rect 5780 3836 6088 3845
rect 5780 3834 5786 3836
rect 5842 3834 5866 3836
rect 5922 3834 5946 3836
rect 6002 3834 6026 3836
rect 6082 3834 6088 3836
rect 5842 3782 5844 3834
rect 6024 3782 6026 3834
rect 5780 3780 5786 3782
rect 5842 3780 5866 3782
rect 5922 3780 5946 3782
rect 6002 3780 6026 3782
rect 6082 3780 6088 3782
rect 5780 3771 6088 3780
rect 7712 3836 8020 3845
rect 7712 3834 7718 3836
rect 7774 3834 7798 3836
rect 7854 3834 7878 3836
rect 7934 3834 7958 3836
rect 8014 3834 8020 3836
rect 7774 3782 7776 3834
rect 7956 3782 7958 3834
rect 7712 3780 7718 3782
rect 7774 3780 7798 3782
rect 7854 3780 7878 3782
rect 7934 3780 7958 3782
rect 8014 3780 8020 3782
rect 7712 3771 8020 3780
rect 2576 3292 2884 3301
rect 2576 3290 2582 3292
rect 2638 3290 2662 3292
rect 2718 3290 2742 3292
rect 2798 3290 2822 3292
rect 2878 3290 2884 3292
rect 2638 3238 2640 3290
rect 2820 3238 2822 3290
rect 2576 3236 2582 3238
rect 2638 3236 2662 3238
rect 2718 3236 2742 3238
rect 2798 3236 2822 3238
rect 2878 3236 2884 3238
rect 2576 3227 2884 3236
rect 4508 3292 4816 3301
rect 4508 3290 4514 3292
rect 4570 3290 4594 3292
rect 4650 3290 4674 3292
rect 4730 3290 4754 3292
rect 4810 3290 4816 3292
rect 4570 3238 4572 3290
rect 4752 3238 4754 3290
rect 4508 3236 4514 3238
rect 4570 3236 4594 3238
rect 4650 3236 4674 3238
rect 4730 3236 4754 3238
rect 4810 3236 4816 3238
rect 4508 3227 4816 3236
rect 6440 3292 6748 3301
rect 6440 3290 6446 3292
rect 6502 3290 6526 3292
rect 6582 3290 6606 3292
rect 6662 3290 6686 3292
rect 6742 3290 6748 3292
rect 6502 3238 6504 3290
rect 6684 3238 6686 3290
rect 6440 3236 6446 3238
rect 6502 3236 6526 3238
rect 6582 3236 6606 3238
rect 6662 3236 6686 3238
rect 6742 3236 6748 3238
rect 6440 3227 6748 3236
rect 8372 3292 8680 3301
rect 8372 3290 8378 3292
rect 8434 3290 8458 3292
rect 8514 3290 8538 3292
rect 8594 3290 8618 3292
rect 8674 3290 8680 3292
rect 8434 3238 8436 3290
rect 8616 3238 8618 3290
rect 8372 3236 8378 3238
rect 8434 3236 8458 3238
rect 8514 3236 8538 3238
rect 8594 3236 8618 3238
rect 8674 3236 8680 3238
rect 8372 3227 8680 3236
rect 1916 2748 2224 2757
rect 1916 2746 1922 2748
rect 1978 2746 2002 2748
rect 2058 2746 2082 2748
rect 2138 2746 2162 2748
rect 2218 2746 2224 2748
rect 1978 2694 1980 2746
rect 2160 2694 2162 2746
rect 1916 2692 1922 2694
rect 1978 2692 2002 2694
rect 2058 2692 2082 2694
rect 2138 2692 2162 2694
rect 2218 2692 2224 2694
rect 1916 2683 2224 2692
rect 3848 2748 4156 2757
rect 3848 2746 3854 2748
rect 3910 2746 3934 2748
rect 3990 2746 4014 2748
rect 4070 2746 4094 2748
rect 4150 2746 4156 2748
rect 3910 2694 3912 2746
rect 4092 2694 4094 2746
rect 3848 2692 3854 2694
rect 3910 2692 3934 2694
rect 3990 2692 4014 2694
rect 4070 2692 4094 2694
rect 4150 2692 4156 2694
rect 3848 2683 4156 2692
rect 5780 2748 6088 2757
rect 5780 2746 5786 2748
rect 5842 2746 5866 2748
rect 5922 2746 5946 2748
rect 6002 2746 6026 2748
rect 6082 2746 6088 2748
rect 5842 2694 5844 2746
rect 6024 2694 6026 2746
rect 5780 2692 5786 2694
rect 5842 2692 5866 2694
rect 5922 2692 5946 2694
rect 6002 2692 6026 2694
rect 6082 2692 6088 2694
rect 5780 2683 6088 2692
rect 7712 2748 8020 2757
rect 7712 2746 7718 2748
rect 7774 2746 7798 2748
rect 7854 2746 7878 2748
rect 7934 2746 7958 2748
rect 8014 2746 8020 2748
rect 7774 2694 7776 2746
rect 7956 2694 7958 2746
rect 7712 2692 7718 2694
rect 7774 2692 7798 2694
rect 7854 2692 7878 2694
rect 7934 2692 7958 2694
rect 8014 2692 8020 2694
rect 7712 2683 8020 2692
rect 2576 2204 2884 2213
rect 2576 2202 2582 2204
rect 2638 2202 2662 2204
rect 2718 2202 2742 2204
rect 2798 2202 2822 2204
rect 2878 2202 2884 2204
rect 2638 2150 2640 2202
rect 2820 2150 2822 2202
rect 2576 2148 2582 2150
rect 2638 2148 2662 2150
rect 2718 2148 2742 2150
rect 2798 2148 2822 2150
rect 2878 2148 2884 2150
rect 2576 2139 2884 2148
rect 4508 2204 4816 2213
rect 4508 2202 4514 2204
rect 4570 2202 4594 2204
rect 4650 2202 4674 2204
rect 4730 2202 4754 2204
rect 4810 2202 4816 2204
rect 4570 2150 4572 2202
rect 4752 2150 4754 2202
rect 4508 2148 4514 2150
rect 4570 2148 4594 2150
rect 4650 2148 4674 2150
rect 4730 2148 4754 2150
rect 4810 2148 4816 2150
rect 4508 2139 4816 2148
rect 6440 2204 6748 2213
rect 6440 2202 6446 2204
rect 6502 2202 6526 2204
rect 6582 2202 6606 2204
rect 6662 2202 6686 2204
rect 6742 2202 6748 2204
rect 6502 2150 6504 2202
rect 6684 2150 6686 2202
rect 6440 2148 6446 2150
rect 6502 2148 6526 2150
rect 6582 2148 6606 2150
rect 6662 2148 6686 2150
rect 6742 2148 6748 2150
rect 6440 2139 6748 2148
rect 8372 2204 8680 2213
rect 8372 2202 8378 2204
rect 8434 2202 8458 2204
rect 8514 2202 8538 2204
rect 8594 2202 8618 2204
rect 8674 2202 8680 2204
rect 8434 2150 8436 2202
rect 8616 2150 8618 2202
rect 8372 2148 8378 2150
rect 8434 2148 8458 2150
rect 8514 2148 8538 2150
rect 8594 2148 8618 2150
rect 8674 2148 8680 2150
rect 8372 2139 8680 2148
<< via2 >>
rect 2582 7642 2638 7644
rect 2662 7642 2718 7644
rect 2742 7642 2798 7644
rect 2822 7642 2878 7644
rect 2582 7590 2628 7642
rect 2628 7590 2638 7642
rect 2662 7590 2692 7642
rect 2692 7590 2704 7642
rect 2704 7590 2718 7642
rect 2742 7590 2756 7642
rect 2756 7590 2768 7642
rect 2768 7590 2798 7642
rect 2822 7590 2832 7642
rect 2832 7590 2878 7642
rect 2582 7588 2638 7590
rect 2662 7588 2718 7590
rect 2742 7588 2798 7590
rect 2822 7588 2878 7590
rect 4514 7642 4570 7644
rect 4594 7642 4650 7644
rect 4674 7642 4730 7644
rect 4754 7642 4810 7644
rect 4514 7590 4560 7642
rect 4560 7590 4570 7642
rect 4594 7590 4624 7642
rect 4624 7590 4636 7642
rect 4636 7590 4650 7642
rect 4674 7590 4688 7642
rect 4688 7590 4700 7642
rect 4700 7590 4730 7642
rect 4754 7590 4764 7642
rect 4764 7590 4810 7642
rect 4514 7588 4570 7590
rect 4594 7588 4650 7590
rect 4674 7588 4730 7590
rect 4754 7588 4810 7590
rect 6446 7642 6502 7644
rect 6526 7642 6582 7644
rect 6606 7642 6662 7644
rect 6686 7642 6742 7644
rect 6446 7590 6492 7642
rect 6492 7590 6502 7642
rect 6526 7590 6556 7642
rect 6556 7590 6568 7642
rect 6568 7590 6582 7642
rect 6606 7590 6620 7642
rect 6620 7590 6632 7642
rect 6632 7590 6662 7642
rect 6686 7590 6696 7642
rect 6696 7590 6742 7642
rect 6446 7588 6502 7590
rect 6526 7588 6582 7590
rect 6606 7588 6662 7590
rect 6686 7588 6742 7590
rect 8378 7642 8434 7644
rect 8458 7642 8514 7644
rect 8538 7642 8594 7644
rect 8618 7642 8674 7644
rect 8378 7590 8424 7642
rect 8424 7590 8434 7642
rect 8458 7590 8488 7642
rect 8488 7590 8500 7642
rect 8500 7590 8514 7642
rect 8538 7590 8552 7642
rect 8552 7590 8564 7642
rect 8564 7590 8594 7642
rect 8618 7590 8628 7642
rect 8628 7590 8674 7642
rect 8378 7588 8434 7590
rect 8458 7588 8514 7590
rect 8538 7588 8594 7590
rect 8618 7588 8674 7590
rect 1922 7098 1978 7100
rect 2002 7098 2058 7100
rect 2082 7098 2138 7100
rect 2162 7098 2218 7100
rect 1922 7046 1968 7098
rect 1968 7046 1978 7098
rect 2002 7046 2032 7098
rect 2032 7046 2044 7098
rect 2044 7046 2058 7098
rect 2082 7046 2096 7098
rect 2096 7046 2108 7098
rect 2108 7046 2138 7098
rect 2162 7046 2172 7098
rect 2172 7046 2218 7098
rect 1922 7044 1978 7046
rect 2002 7044 2058 7046
rect 2082 7044 2138 7046
rect 2162 7044 2218 7046
rect 3854 7098 3910 7100
rect 3934 7098 3990 7100
rect 4014 7098 4070 7100
rect 4094 7098 4150 7100
rect 3854 7046 3900 7098
rect 3900 7046 3910 7098
rect 3934 7046 3964 7098
rect 3964 7046 3976 7098
rect 3976 7046 3990 7098
rect 4014 7046 4028 7098
rect 4028 7046 4040 7098
rect 4040 7046 4070 7098
rect 4094 7046 4104 7098
rect 4104 7046 4150 7098
rect 3854 7044 3910 7046
rect 3934 7044 3990 7046
rect 4014 7044 4070 7046
rect 4094 7044 4150 7046
rect 5786 7098 5842 7100
rect 5866 7098 5922 7100
rect 5946 7098 6002 7100
rect 6026 7098 6082 7100
rect 5786 7046 5832 7098
rect 5832 7046 5842 7098
rect 5866 7046 5896 7098
rect 5896 7046 5908 7098
rect 5908 7046 5922 7098
rect 5946 7046 5960 7098
rect 5960 7046 5972 7098
rect 5972 7046 6002 7098
rect 6026 7046 6036 7098
rect 6036 7046 6082 7098
rect 5786 7044 5842 7046
rect 5866 7044 5922 7046
rect 5946 7044 6002 7046
rect 6026 7044 6082 7046
rect 7718 7098 7774 7100
rect 7798 7098 7854 7100
rect 7878 7098 7934 7100
rect 7958 7098 8014 7100
rect 7718 7046 7764 7098
rect 7764 7046 7774 7098
rect 7798 7046 7828 7098
rect 7828 7046 7840 7098
rect 7840 7046 7854 7098
rect 7878 7046 7892 7098
rect 7892 7046 7904 7098
rect 7904 7046 7934 7098
rect 7958 7046 7968 7098
rect 7968 7046 8014 7098
rect 7718 7044 7774 7046
rect 7798 7044 7854 7046
rect 7878 7044 7934 7046
rect 7958 7044 8014 7046
rect 2582 6554 2638 6556
rect 2662 6554 2718 6556
rect 2742 6554 2798 6556
rect 2822 6554 2878 6556
rect 2582 6502 2628 6554
rect 2628 6502 2638 6554
rect 2662 6502 2692 6554
rect 2692 6502 2704 6554
rect 2704 6502 2718 6554
rect 2742 6502 2756 6554
rect 2756 6502 2768 6554
rect 2768 6502 2798 6554
rect 2822 6502 2832 6554
rect 2832 6502 2878 6554
rect 2582 6500 2638 6502
rect 2662 6500 2718 6502
rect 2742 6500 2798 6502
rect 2822 6500 2878 6502
rect 4514 6554 4570 6556
rect 4594 6554 4650 6556
rect 4674 6554 4730 6556
rect 4754 6554 4810 6556
rect 4514 6502 4560 6554
rect 4560 6502 4570 6554
rect 4594 6502 4624 6554
rect 4624 6502 4636 6554
rect 4636 6502 4650 6554
rect 4674 6502 4688 6554
rect 4688 6502 4700 6554
rect 4700 6502 4730 6554
rect 4754 6502 4764 6554
rect 4764 6502 4810 6554
rect 4514 6500 4570 6502
rect 4594 6500 4650 6502
rect 4674 6500 4730 6502
rect 4754 6500 4810 6502
rect 6446 6554 6502 6556
rect 6526 6554 6582 6556
rect 6606 6554 6662 6556
rect 6686 6554 6742 6556
rect 6446 6502 6492 6554
rect 6492 6502 6502 6554
rect 6526 6502 6556 6554
rect 6556 6502 6568 6554
rect 6568 6502 6582 6554
rect 6606 6502 6620 6554
rect 6620 6502 6632 6554
rect 6632 6502 6662 6554
rect 6686 6502 6696 6554
rect 6696 6502 6742 6554
rect 6446 6500 6502 6502
rect 6526 6500 6582 6502
rect 6606 6500 6662 6502
rect 6686 6500 6742 6502
rect 8378 6554 8434 6556
rect 8458 6554 8514 6556
rect 8538 6554 8594 6556
rect 8618 6554 8674 6556
rect 8378 6502 8424 6554
rect 8424 6502 8434 6554
rect 8458 6502 8488 6554
rect 8488 6502 8500 6554
rect 8500 6502 8514 6554
rect 8538 6502 8552 6554
rect 8552 6502 8564 6554
rect 8564 6502 8594 6554
rect 8618 6502 8628 6554
rect 8628 6502 8674 6554
rect 8378 6500 8434 6502
rect 8458 6500 8514 6502
rect 8538 6500 8594 6502
rect 8618 6500 8674 6502
rect 1922 6010 1978 6012
rect 2002 6010 2058 6012
rect 2082 6010 2138 6012
rect 2162 6010 2218 6012
rect 1922 5958 1968 6010
rect 1968 5958 1978 6010
rect 2002 5958 2032 6010
rect 2032 5958 2044 6010
rect 2044 5958 2058 6010
rect 2082 5958 2096 6010
rect 2096 5958 2108 6010
rect 2108 5958 2138 6010
rect 2162 5958 2172 6010
rect 2172 5958 2218 6010
rect 1922 5956 1978 5958
rect 2002 5956 2058 5958
rect 2082 5956 2138 5958
rect 2162 5956 2218 5958
rect 3854 6010 3910 6012
rect 3934 6010 3990 6012
rect 4014 6010 4070 6012
rect 4094 6010 4150 6012
rect 3854 5958 3900 6010
rect 3900 5958 3910 6010
rect 3934 5958 3964 6010
rect 3964 5958 3976 6010
rect 3976 5958 3990 6010
rect 4014 5958 4028 6010
rect 4028 5958 4040 6010
rect 4040 5958 4070 6010
rect 4094 5958 4104 6010
rect 4104 5958 4150 6010
rect 3854 5956 3910 5958
rect 3934 5956 3990 5958
rect 4014 5956 4070 5958
rect 4094 5956 4150 5958
rect 5786 6010 5842 6012
rect 5866 6010 5922 6012
rect 5946 6010 6002 6012
rect 6026 6010 6082 6012
rect 5786 5958 5832 6010
rect 5832 5958 5842 6010
rect 5866 5958 5896 6010
rect 5896 5958 5908 6010
rect 5908 5958 5922 6010
rect 5946 5958 5960 6010
rect 5960 5958 5972 6010
rect 5972 5958 6002 6010
rect 6026 5958 6036 6010
rect 6036 5958 6082 6010
rect 5786 5956 5842 5958
rect 5866 5956 5922 5958
rect 5946 5956 6002 5958
rect 6026 5956 6082 5958
rect 7718 6010 7774 6012
rect 7798 6010 7854 6012
rect 7878 6010 7934 6012
rect 7958 6010 8014 6012
rect 7718 5958 7764 6010
rect 7764 5958 7774 6010
rect 7798 5958 7828 6010
rect 7828 5958 7840 6010
rect 7840 5958 7854 6010
rect 7878 5958 7892 6010
rect 7892 5958 7904 6010
rect 7904 5958 7934 6010
rect 7958 5958 7968 6010
rect 7968 5958 8014 6010
rect 7718 5956 7774 5958
rect 7798 5956 7854 5958
rect 7878 5956 7934 5958
rect 7958 5956 8014 5958
rect 1398 5480 1454 5536
rect 2582 5466 2638 5468
rect 2662 5466 2718 5468
rect 2742 5466 2798 5468
rect 2822 5466 2878 5468
rect 2582 5414 2628 5466
rect 2628 5414 2638 5466
rect 2662 5414 2692 5466
rect 2692 5414 2704 5466
rect 2704 5414 2718 5466
rect 2742 5414 2756 5466
rect 2756 5414 2768 5466
rect 2768 5414 2798 5466
rect 2822 5414 2832 5466
rect 2832 5414 2878 5466
rect 2582 5412 2638 5414
rect 2662 5412 2718 5414
rect 2742 5412 2798 5414
rect 2822 5412 2878 5414
rect 1922 4922 1978 4924
rect 2002 4922 2058 4924
rect 2082 4922 2138 4924
rect 2162 4922 2218 4924
rect 1922 4870 1968 4922
rect 1968 4870 1978 4922
rect 2002 4870 2032 4922
rect 2032 4870 2044 4922
rect 2044 4870 2058 4922
rect 2082 4870 2096 4922
rect 2096 4870 2108 4922
rect 2108 4870 2138 4922
rect 2162 4870 2172 4922
rect 2172 4870 2218 4922
rect 1922 4868 1978 4870
rect 2002 4868 2058 4870
rect 2082 4868 2138 4870
rect 2162 4868 2218 4870
rect 3854 4922 3910 4924
rect 3934 4922 3990 4924
rect 4014 4922 4070 4924
rect 4094 4922 4150 4924
rect 3854 4870 3900 4922
rect 3900 4870 3910 4922
rect 3934 4870 3964 4922
rect 3964 4870 3976 4922
rect 3976 4870 3990 4922
rect 4014 4870 4028 4922
rect 4028 4870 4040 4922
rect 4040 4870 4070 4922
rect 4094 4870 4104 4922
rect 4104 4870 4150 4922
rect 3854 4868 3910 4870
rect 3934 4868 3990 4870
rect 4014 4868 4070 4870
rect 4094 4868 4150 4870
rect 938 4800 994 4856
rect 4514 5466 4570 5468
rect 4594 5466 4650 5468
rect 4674 5466 4730 5468
rect 4754 5466 4810 5468
rect 4514 5414 4560 5466
rect 4560 5414 4570 5466
rect 4594 5414 4624 5466
rect 4624 5414 4636 5466
rect 4636 5414 4650 5466
rect 4674 5414 4688 5466
rect 4688 5414 4700 5466
rect 4700 5414 4730 5466
rect 4754 5414 4764 5466
rect 4764 5414 4810 5466
rect 4514 5412 4570 5414
rect 4594 5412 4650 5414
rect 4674 5412 4730 5414
rect 4754 5412 4810 5414
rect 6446 5466 6502 5468
rect 6526 5466 6582 5468
rect 6606 5466 6662 5468
rect 6686 5466 6742 5468
rect 6446 5414 6492 5466
rect 6492 5414 6502 5466
rect 6526 5414 6556 5466
rect 6556 5414 6568 5466
rect 6568 5414 6582 5466
rect 6606 5414 6620 5466
rect 6620 5414 6632 5466
rect 6632 5414 6662 5466
rect 6686 5414 6696 5466
rect 6696 5414 6742 5466
rect 6446 5412 6502 5414
rect 6526 5412 6582 5414
rect 6606 5412 6662 5414
rect 6686 5412 6742 5414
rect 8758 5516 8760 5536
rect 8760 5516 8812 5536
rect 8812 5516 8814 5536
rect 8758 5480 8814 5516
rect 8378 5466 8434 5468
rect 8458 5466 8514 5468
rect 8538 5466 8594 5468
rect 8618 5466 8674 5468
rect 8378 5414 8424 5466
rect 8424 5414 8434 5466
rect 8458 5414 8488 5466
rect 8488 5414 8500 5466
rect 8500 5414 8514 5466
rect 8538 5414 8552 5466
rect 8552 5414 8564 5466
rect 8564 5414 8594 5466
rect 8618 5414 8628 5466
rect 8628 5414 8674 5466
rect 8378 5412 8434 5414
rect 8458 5412 8514 5414
rect 8538 5412 8594 5414
rect 8618 5412 8674 5414
rect 5786 4922 5842 4924
rect 5866 4922 5922 4924
rect 5946 4922 6002 4924
rect 6026 4922 6082 4924
rect 5786 4870 5832 4922
rect 5832 4870 5842 4922
rect 5866 4870 5896 4922
rect 5896 4870 5908 4922
rect 5908 4870 5922 4922
rect 5946 4870 5960 4922
rect 5960 4870 5972 4922
rect 5972 4870 6002 4922
rect 6026 4870 6036 4922
rect 6036 4870 6082 4922
rect 5786 4868 5842 4870
rect 5866 4868 5922 4870
rect 5946 4868 6002 4870
rect 6026 4868 6082 4870
rect 7718 4922 7774 4924
rect 7798 4922 7854 4924
rect 7878 4922 7934 4924
rect 7958 4922 8014 4924
rect 7718 4870 7764 4922
rect 7764 4870 7774 4922
rect 7798 4870 7828 4922
rect 7828 4870 7840 4922
rect 7840 4870 7854 4922
rect 7878 4870 7892 4922
rect 7892 4870 7904 4922
rect 7904 4870 7934 4922
rect 7958 4870 7968 4922
rect 7968 4870 8014 4922
rect 7718 4868 7774 4870
rect 7798 4868 7854 4870
rect 7878 4868 7934 4870
rect 7958 4868 8014 4870
rect 8390 4800 8446 4856
rect 2582 4378 2638 4380
rect 2662 4378 2718 4380
rect 2742 4378 2798 4380
rect 2822 4378 2878 4380
rect 2582 4326 2628 4378
rect 2628 4326 2638 4378
rect 2662 4326 2692 4378
rect 2692 4326 2704 4378
rect 2704 4326 2718 4378
rect 2742 4326 2756 4378
rect 2756 4326 2768 4378
rect 2768 4326 2798 4378
rect 2822 4326 2832 4378
rect 2832 4326 2878 4378
rect 2582 4324 2638 4326
rect 2662 4324 2718 4326
rect 2742 4324 2798 4326
rect 2822 4324 2878 4326
rect 4514 4378 4570 4380
rect 4594 4378 4650 4380
rect 4674 4378 4730 4380
rect 4754 4378 4810 4380
rect 4514 4326 4560 4378
rect 4560 4326 4570 4378
rect 4594 4326 4624 4378
rect 4624 4326 4636 4378
rect 4636 4326 4650 4378
rect 4674 4326 4688 4378
rect 4688 4326 4700 4378
rect 4700 4326 4730 4378
rect 4754 4326 4764 4378
rect 4764 4326 4810 4378
rect 4514 4324 4570 4326
rect 4594 4324 4650 4326
rect 4674 4324 4730 4326
rect 4754 4324 4810 4326
rect 6446 4378 6502 4380
rect 6526 4378 6582 4380
rect 6606 4378 6662 4380
rect 6686 4378 6742 4380
rect 6446 4326 6492 4378
rect 6492 4326 6502 4378
rect 6526 4326 6556 4378
rect 6556 4326 6568 4378
rect 6568 4326 6582 4378
rect 6606 4326 6620 4378
rect 6620 4326 6632 4378
rect 6632 4326 6662 4378
rect 6686 4326 6696 4378
rect 6696 4326 6742 4378
rect 6446 4324 6502 4326
rect 6526 4324 6582 4326
rect 6606 4324 6662 4326
rect 6686 4324 6742 4326
rect 8378 4378 8434 4380
rect 8458 4378 8514 4380
rect 8538 4378 8594 4380
rect 8618 4378 8674 4380
rect 8378 4326 8424 4378
rect 8424 4326 8434 4378
rect 8458 4326 8488 4378
rect 8488 4326 8500 4378
rect 8500 4326 8514 4378
rect 8538 4326 8552 4378
rect 8552 4326 8564 4378
rect 8564 4326 8594 4378
rect 8618 4326 8628 4378
rect 8628 4326 8674 4378
rect 8378 4324 8434 4326
rect 8458 4324 8514 4326
rect 8538 4324 8594 4326
rect 8618 4324 8674 4326
rect 938 4120 994 4176
rect 1922 3834 1978 3836
rect 2002 3834 2058 3836
rect 2082 3834 2138 3836
rect 2162 3834 2218 3836
rect 1922 3782 1968 3834
rect 1968 3782 1978 3834
rect 2002 3782 2032 3834
rect 2032 3782 2044 3834
rect 2044 3782 2058 3834
rect 2082 3782 2096 3834
rect 2096 3782 2108 3834
rect 2108 3782 2138 3834
rect 2162 3782 2172 3834
rect 2172 3782 2218 3834
rect 1922 3780 1978 3782
rect 2002 3780 2058 3782
rect 2082 3780 2138 3782
rect 2162 3780 2218 3782
rect 3854 3834 3910 3836
rect 3934 3834 3990 3836
rect 4014 3834 4070 3836
rect 4094 3834 4150 3836
rect 3854 3782 3900 3834
rect 3900 3782 3910 3834
rect 3934 3782 3964 3834
rect 3964 3782 3976 3834
rect 3976 3782 3990 3834
rect 4014 3782 4028 3834
rect 4028 3782 4040 3834
rect 4040 3782 4070 3834
rect 4094 3782 4104 3834
rect 4104 3782 4150 3834
rect 3854 3780 3910 3782
rect 3934 3780 3990 3782
rect 4014 3780 4070 3782
rect 4094 3780 4150 3782
rect 5786 3834 5842 3836
rect 5866 3834 5922 3836
rect 5946 3834 6002 3836
rect 6026 3834 6082 3836
rect 5786 3782 5832 3834
rect 5832 3782 5842 3834
rect 5866 3782 5896 3834
rect 5896 3782 5908 3834
rect 5908 3782 5922 3834
rect 5946 3782 5960 3834
rect 5960 3782 5972 3834
rect 5972 3782 6002 3834
rect 6026 3782 6036 3834
rect 6036 3782 6082 3834
rect 5786 3780 5842 3782
rect 5866 3780 5922 3782
rect 5946 3780 6002 3782
rect 6026 3780 6082 3782
rect 7718 3834 7774 3836
rect 7798 3834 7854 3836
rect 7878 3834 7934 3836
rect 7958 3834 8014 3836
rect 7718 3782 7764 3834
rect 7764 3782 7774 3834
rect 7798 3782 7828 3834
rect 7828 3782 7840 3834
rect 7840 3782 7854 3834
rect 7878 3782 7892 3834
rect 7892 3782 7904 3834
rect 7904 3782 7934 3834
rect 7958 3782 7968 3834
rect 7968 3782 8014 3834
rect 7718 3780 7774 3782
rect 7798 3780 7854 3782
rect 7878 3780 7934 3782
rect 7958 3780 8014 3782
rect 2582 3290 2638 3292
rect 2662 3290 2718 3292
rect 2742 3290 2798 3292
rect 2822 3290 2878 3292
rect 2582 3238 2628 3290
rect 2628 3238 2638 3290
rect 2662 3238 2692 3290
rect 2692 3238 2704 3290
rect 2704 3238 2718 3290
rect 2742 3238 2756 3290
rect 2756 3238 2768 3290
rect 2768 3238 2798 3290
rect 2822 3238 2832 3290
rect 2832 3238 2878 3290
rect 2582 3236 2638 3238
rect 2662 3236 2718 3238
rect 2742 3236 2798 3238
rect 2822 3236 2878 3238
rect 4514 3290 4570 3292
rect 4594 3290 4650 3292
rect 4674 3290 4730 3292
rect 4754 3290 4810 3292
rect 4514 3238 4560 3290
rect 4560 3238 4570 3290
rect 4594 3238 4624 3290
rect 4624 3238 4636 3290
rect 4636 3238 4650 3290
rect 4674 3238 4688 3290
rect 4688 3238 4700 3290
rect 4700 3238 4730 3290
rect 4754 3238 4764 3290
rect 4764 3238 4810 3290
rect 4514 3236 4570 3238
rect 4594 3236 4650 3238
rect 4674 3236 4730 3238
rect 4754 3236 4810 3238
rect 6446 3290 6502 3292
rect 6526 3290 6582 3292
rect 6606 3290 6662 3292
rect 6686 3290 6742 3292
rect 6446 3238 6492 3290
rect 6492 3238 6502 3290
rect 6526 3238 6556 3290
rect 6556 3238 6568 3290
rect 6568 3238 6582 3290
rect 6606 3238 6620 3290
rect 6620 3238 6632 3290
rect 6632 3238 6662 3290
rect 6686 3238 6696 3290
rect 6696 3238 6742 3290
rect 6446 3236 6502 3238
rect 6526 3236 6582 3238
rect 6606 3236 6662 3238
rect 6686 3236 6742 3238
rect 8378 3290 8434 3292
rect 8458 3290 8514 3292
rect 8538 3290 8594 3292
rect 8618 3290 8674 3292
rect 8378 3238 8424 3290
rect 8424 3238 8434 3290
rect 8458 3238 8488 3290
rect 8488 3238 8500 3290
rect 8500 3238 8514 3290
rect 8538 3238 8552 3290
rect 8552 3238 8564 3290
rect 8564 3238 8594 3290
rect 8618 3238 8628 3290
rect 8628 3238 8674 3290
rect 8378 3236 8434 3238
rect 8458 3236 8514 3238
rect 8538 3236 8594 3238
rect 8618 3236 8674 3238
rect 1922 2746 1978 2748
rect 2002 2746 2058 2748
rect 2082 2746 2138 2748
rect 2162 2746 2218 2748
rect 1922 2694 1968 2746
rect 1968 2694 1978 2746
rect 2002 2694 2032 2746
rect 2032 2694 2044 2746
rect 2044 2694 2058 2746
rect 2082 2694 2096 2746
rect 2096 2694 2108 2746
rect 2108 2694 2138 2746
rect 2162 2694 2172 2746
rect 2172 2694 2218 2746
rect 1922 2692 1978 2694
rect 2002 2692 2058 2694
rect 2082 2692 2138 2694
rect 2162 2692 2218 2694
rect 3854 2746 3910 2748
rect 3934 2746 3990 2748
rect 4014 2746 4070 2748
rect 4094 2746 4150 2748
rect 3854 2694 3900 2746
rect 3900 2694 3910 2746
rect 3934 2694 3964 2746
rect 3964 2694 3976 2746
rect 3976 2694 3990 2746
rect 4014 2694 4028 2746
rect 4028 2694 4040 2746
rect 4040 2694 4070 2746
rect 4094 2694 4104 2746
rect 4104 2694 4150 2746
rect 3854 2692 3910 2694
rect 3934 2692 3990 2694
rect 4014 2692 4070 2694
rect 4094 2692 4150 2694
rect 5786 2746 5842 2748
rect 5866 2746 5922 2748
rect 5946 2746 6002 2748
rect 6026 2746 6082 2748
rect 5786 2694 5832 2746
rect 5832 2694 5842 2746
rect 5866 2694 5896 2746
rect 5896 2694 5908 2746
rect 5908 2694 5922 2746
rect 5946 2694 5960 2746
rect 5960 2694 5972 2746
rect 5972 2694 6002 2746
rect 6026 2694 6036 2746
rect 6036 2694 6082 2746
rect 5786 2692 5842 2694
rect 5866 2692 5922 2694
rect 5946 2692 6002 2694
rect 6026 2692 6082 2694
rect 7718 2746 7774 2748
rect 7798 2746 7854 2748
rect 7878 2746 7934 2748
rect 7958 2746 8014 2748
rect 7718 2694 7764 2746
rect 7764 2694 7774 2746
rect 7798 2694 7828 2746
rect 7828 2694 7840 2746
rect 7840 2694 7854 2746
rect 7878 2694 7892 2746
rect 7892 2694 7904 2746
rect 7904 2694 7934 2746
rect 7958 2694 7968 2746
rect 7968 2694 8014 2746
rect 7718 2692 7774 2694
rect 7798 2692 7854 2694
rect 7878 2692 7934 2694
rect 7958 2692 8014 2694
rect 2582 2202 2638 2204
rect 2662 2202 2718 2204
rect 2742 2202 2798 2204
rect 2822 2202 2878 2204
rect 2582 2150 2628 2202
rect 2628 2150 2638 2202
rect 2662 2150 2692 2202
rect 2692 2150 2704 2202
rect 2704 2150 2718 2202
rect 2742 2150 2756 2202
rect 2756 2150 2768 2202
rect 2768 2150 2798 2202
rect 2822 2150 2832 2202
rect 2832 2150 2878 2202
rect 2582 2148 2638 2150
rect 2662 2148 2718 2150
rect 2742 2148 2798 2150
rect 2822 2148 2878 2150
rect 4514 2202 4570 2204
rect 4594 2202 4650 2204
rect 4674 2202 4730 2204
rect 4754 2202 4810 2204
rect 4514 2150 4560 2202
rect 4560 2150 4570 2202
rect 4594 2150 4624 2202
rect 4624 2150 4636 2202
rect 4636 2150 4650 2202
rect 4674 2150 4688 2202
rect 4688 2150 4700 2202
rect 4700 2150 4730 2202
rect 4754 2150 4764 2202
rect 4764 2150 4810 2202
rect 4514 2148 4570 2150
rect 4594 2148 4650 2150
rect 4674 2148 4730 2150
rect 4754 2148 4810 2150
rect 6446 2202 6502 2204
rect 6526 2202 6582 2204
rect 6606 2202 6662 2204
rect 6686 2202 6742 2204
rect 6446 2150 6492 2202
rect 6492 2150 6502 2202
rect 6526 2150 6556 2202
rect 6556 2150 6568 2202
rect 6568 2150 6582 2202
rect 6606 2150 6620 2202
rect 6620 2150 6632 2202
rect 6632 2150 6662 2202
rect 6686 2150 6696 2202
rect 6696 2150 6742 2202
rect 6446 2148 6502 2150
rect 6526 2148 6582 2150
rect 6606 2148 6662 2150
rect 6686 2148 6742 2150
rect 8378 2202 8434 2204
rect 8458 2202 8514 2204
rect 8538 2202 8594 2204
rect 8618 2202 8674 2204
rect 8378 2150 8424 2202
rect 8424 2150 8434 2202
rect 8458 2150 8488 2202
rect 8488 2150 8500 2202
rect 8500 2150 8514 2202
rect 8538 2150 8552 2202
rect 8552 2150 8564 2202
rect 8564 2150 8594 2202
rect 8618 2150 8628 2202
rect 8628 2150 8674 2202
rect 8378 2148 8434 2150
rect 8458 2148 8514 2150
rect 8538 2148 8594 2150
rect 8618 2148 8674 2150
<< metal3 >>
rect 2572 7648 2888 7649
rect 2572 7584 2578 7648
rect 2642 7584 2658 7648
rect 2722 7584 2738 7648
rect 2802 7584 2818 7648
rect 2882 7584 2888 7648
rect 2572 7583 2888 7584
rect 4504 7648 4820 7649
rect 4504 7584 4510 7648
rect 4574 7584 4590 7648
rect 4654 7584 4670 7648
rect 4734 7584 4750 7648
rect 4814 7584 4820 7648
rect 4504 7583 4820 7584
rect 6436 7648 6752 7649
rect 6436 7584 6442 7648
rect 6506 7584 6522 7648
rect 6586 7584 6602 7648
rect 6666 7584 6682 7648
rect 6746 7584 6752 7648
rect 6436 7583 6752 7584
rect 8368 7648 8684 7649
rect 8368 7584 8374 7648
rect 8438 7584 8454 7648
rect 8518 7584 8534 7648
rect 8598 7584 8614 7648
rect 8678 7584 8684 7648
rect 8368 7583 8684 7584
rect 1912 7104 2228 7105
rect 1912 7040 1918 7104
rect 1982 7040 1998 7104
rect 2062 7040 2078 7104
rect 2142 7040 2158 7104
rect 2222 7040 2228 7104
rect 1912 7039 2228 7040
rect 3844 7104 4160 7105
rect 3844 7040 3850 7104
rect 3914 7040 3930 7104
rect 3994 7040 4010 7104
rect 4074 7040 4090 7104
rect 4154 7040 4160 7104
rect 3844 7039 4160 7040
rect 5776 7104 6092 7105
rect 5776 7040 5782 7104
rect 5846 7040 5862 7104
rect 5926 7040 5942 7104
rect 6006 7040 6022 7104
rect 6086 7040 6092 7104
rect 5776 7039 6092 7040
rect 7708 7104 8024 7105
rect 7708 7040 7714 7104
rect 7778 7040 7794 7104
rect 7858 7040 7874 7104
rect 7938 7040 7954 7104
rect 8018 7040 8024 7104
rect 7708 7039 8024 7040
rect 2572 6560 2888 6561
rect 2572 6496 2578 6560
rect 2642 6496 2658 6560
rect 2722 6496 2738 6560
rect 2802 6496 2818 6560
rect 2882 6496 2888 6560
rect 2572 6495 2888 6496
rect 4504 6560 4820 6561
rect 4504 6496 4510 6560
rect 4574 6496 4590 6560
rect 4654 6496 4670 6560
rect 4734 6496 4750 6560
rect 4814 6496 4820 6560
rect 4504 6495 4820 6496
rect 6436 6560 6752 6561
rect 6436 6496 6442 6560
rect 6506 6496 6522 6560
rect 6586 6496 6602 6560
rect 6666 6496 6682 6560
rect 6746 6496 6752 6560
rect 6436 6495 6752 6496
rect 8368 6560 8684 6561
rect 8368 6496 8374 6560
rect 8438 6496 8454 6560
rect 8518 6496 8534 6560
rect 8598 6496 8614 6560
rect 8678 6496 8684 6560
rect 8368 6495 8684 6496
rect 1912 6016 2228 6017
rect 1912 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2228 6016
rect 1912 5951 2228 5952
rect 3844 6016 4160 6017
rect 3844 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4160 6016
rect 3844 5951 4160 5952
rect 5776 6016 6092 6017
rect 5776 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6092 6016
rect 5776 5951 6092 5952
rect 7708 6016 8024 6017
rect 7708 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8024 6016
rect 7708 5951 8024 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 8753 5538 8819 5541
rect 9200 5538 10000 5568
rect 8753 5536 10000 5538
rect 8753 5480 8758 5536
rect 8814 5480 10000 5536
rect 8753 5478 10000 5480
rect 8753 5475 8819 5478
rect 2572 5472 2888 5473
rect 2572 5408 2578 5472
rect 2642 5408 2658 5472
rect 2722 5408 2738 5472
rect 2802 5408 2818 5472
rect 2882 5408 2888 5472
rect 2572 5407 2888 5408
rect 4504 5472 4820 5473
rect 4504 5408 4510 5472
rect 4574 5408 4590 5472
rect 4654 5408 4670 5472
rect 4734 5408 4750 5472
rect 4814 5408 4820 5472
rect 4504 5407 4820 5408
rect 6436 5472 6752 5473
rect 6436 5408 6442 5472
rect 6506 5408 6522 5472
rect 6586 5408 6602 5472
rect 6666 5408 6682 5472
rect 6746 5408 6752 5472
rect 6436 5407 6752 5408
rect 8368 5472 8684 5473
rect 8368 5408 8374 5472
rect 8438 5408 8454 5472
rect 8518 5408 8534 5472
rect 8598 5408 8614 5472
rect 8678 5408 8684 5472
rect 9200 5448 10000 5478
rect 8368 5407 8684 5408
rect 1912 4928 2228 4929
rect 0 4858 800 4888
rect 1912 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2228 4928
rect 1912 4863 2228 4864
rect 3844 4928 4160 4929
rect 3844 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4160 4928
rect 3844 4863 4160 4864
rect 5776 4928 6092 4929
rect 5776 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6092 4928
rect 5776 4863 6092 4864
rect 7708 4928 8024 4929
rect 7708 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8024 4928
rect 7708 4863 8024 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 8385 4858 8451 4861
rect 9200 4858 10000 4888
rect 8385 4856 10000 4858
rect 8385 4800 8390 4856
rect 8446 4800 10000 4856
rect 8385 4798 10000 4800
rect 8385 4795 8451 4798
rect 9200 4768 10000 4798
rect 2572 4384 2888 4385
rect 2572 4320 2578 4384
rect 2642 4320 2658 4384
rect 2722 4320 2738 4384
rect 2802 4320 2818 4384
rect 2882 4320 2888 4384
rect 2572 4319 2888 4320
rect 4504 4384 4820 4385
rect 4504 4320 4510 4384
rect 4574 4320 4590 4384
rect 4654 4320 4670 4384
rect 4734 4320 4750 4384
rect 4814 4320 4820 4384
rect 4504 4319 4820 4320
rect 6436 4384 6752 4385
rect 6436 4320 6442 4384
rect 6506 4320 6522 4384
rect 6586 4320 6602 4384
rect 6666 4320 6682 4384
rect 6746 4320 6752 4384
rect 6436 4319 6752 4320
rect 8368 4384 8684 4385
rect 8368 4320 8374 4384
rect 8438 4320 8454 4384
rect 8518 4320 8534 4384
rect 8598 4320 8614 4384
rect 8678 4320 8684 4384
rect 8368 4319 8684 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 1912 3840 2228 3841
rect 1912 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2228 3840
rect 1912 3775 2228 3776
rect 3844 3840 4160 3841
rect 3844 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4160 3840
rect 3844 3775 4160 3776
rect 5776 3840 6092 3841
rect 5776 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6092 3840
rect 5776 3775 6092 3776
rect 7708 3840 8024 3841
rect 7708 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8024 3840
rect 7708 3775 8024 3776
rect 2572 3296 2888 3297
rect 2572 3232 2578 3296
rect 2642 3232 2658 3296
rect 2722 3232 2738 3296
rect 2802 3232 2818 3296
rect 2882 3232 2888 3296
rect 2572 3231 2888 3232
rect 4504 3296 4820 3297
rect 4504 3232 4510 3296
rect 4574 3232 4590 3296
rect 4654 3232 4670 3296
rect 4734 3232 4750 3296
rect 4814 3232 4820 3296
rect 4504 3231 4820 3232
rect 6436 3296 6752 3297
rect 6436 3232 6442 3296
rect 6506 3232 6522 3296
rect 6586 3232 6602 3296
rect 6666 3232 6682 3296
rect 6746 3232 6752 3296
rect 6436 3231 6752 3232
rect 8368 3296 8684 3297
rect 8368 3232 8374 3296
rect 8438 3232 8454 3296
rect 8518 3232 8534 3296
rect 8598 3232 8614 3296
rect 8678 3232 8684 3296
rect 8368 3231 8684 3232
rect 1912 2752 2228 2753
rect 1912 2688 1918 2752
rect 1982 2688 1998 2752
rect 2062 2688 2078 2752
rect 2142 2688 2158 2752
rect 2222 2688 2228 2752
rect 1912 2687 2228 2688
rect 3844 2752 4160 2753
rect 3844 2688 3850 2752
rect 3914 2688 3930 2752
rect 3994 2688 4010 2752
rect 4074 2688 4090 2752
rect 4154 2688 4160 2752
rect 3844 2687 4160 2688
rect 5776 2752 6092 2753
rect 5776 2688 5782 2752
rect 5846 2688 5862 2752
rect 5926 2688 5942 2752
rect 6006 2688 6022 2752
rect 6086 2688 6092 2752
rect 5776 2687 6092 2688
rect 7708 2752 8024 2753
rect 7708 2688 7714 2752
rect 7778 2688 7794 2752
rect 7858 2688 7874 2752
rect 7938 2688 7954 2752
rect 8018 2688 8024 2752
rect 7708 2687 8024 2688
rect 2572 2208 2888 2209
rect 2572 2144 2578 2208
rect 2642 2144 2658 2208
rect 2722 2144 2738 2208
rect 2802 2144 2818 2208
rect 2882 2144 2888 2208
rect 2572 2143 2888 2144
rect 4504 2208 4820 2209
rect 4504 2144 4510 2208
rect 4574 2144 4590 2208
rect 4654 2144 4670 2208
rect 4734 2144 4750 2208
rect 4814 2144 4820 2208
rect 4504 2143 4820 2144
rect 6436 2208 6752 2209
rect 6436 2144 6442 2208
rect 6506 2144 6522 2208
rect 6586 2144 6602 2208
rect 6666 2144 6682 2208
rect 6746 2144 6752 2208
rect 6436 2143 6752 2144
rect 8368 2208 8684 2209
rect 8368 2144 8374 2208
rect 8438 2144 8454 2208
rect 8518 2144 8534 2208
rect 8598 2144 8614 2208
rect 8678 2144 8684 2208
rect 8368 2143 8684 2144
<< via3 >>
rect 2578 7644 2642 7648
rect 2578 7588 2582 7644
rect 2582 7588 2638 7644
rect 2638 7588 2642 7644
rect 2578 7584 2642 7588
rect 2658 7644 2722 7648
rect 2658 7588 2662 7644
rect 2662 7588 2718 7644
rect 2718 7588 2722 7644
rect 2658 7584 2722 7588
rect 2738 7644 2802 7648
rect 2738 7588 2742 7644
rect 2742 7588 2798 7644
rect 2798 7588 2802 7644
rect 2738 7584 2802 7588
rect 2818 7644 2882 7648
rect 2818 7588 2822 7644
rect 2822 7588 2878 7644
rect 2878 7588 2882 7644
rect 2818 7584 2882 7588
rect 4510 7644 4574 7648
rect 4510 7588 4514 7644
rect 4514 7588 4570 7644
rect 4570 7588 4574 7644
rect 4510 7584 4574 7588
rect 4590 7644 4654 7648
rect 4590 7588 4594 7644
rect 4594 7588 4650 7644
rect 4650 7588 4654 7644
rect 4590 7584 4654 7588
rect 4670 7644 4734 7648
rect 4670 7588 4674 7644
rect 4674 7588 4730 7644
rect 4730 7588 4734 7644
rect 4670 7584 4734 7588
rect 4750 7644 4814 7648
rect 4750 7588 4754 7644
rect 4754 7588 4810 7644
rect 4810 7588 4814 7644
rect 4750 7584 4814 7588
rect 6442 7644 6506 7648
rect 6442 7588 6446 7644
rect 6446 7588 6502 7644
rect 6502 7588 6506 7644
rect 6442 7584 6506 7588
rect 6522 7644 6586 7648
rect 6522 7588 6526 7644
rect 6526 7588 6582 7644
rect 6582 7588 6586 7644
rect 6522 7584 6586 7588
rect 6602 7644 6666 7648
rect 6602 7588 6606 7644
rect 6606 7588 6662 7644
rect 6662 7588 6666 7644
rect 6602 7584 6666 7588
rect 6682 7644 6746 7648
rect 6682 7588 6686 7644
rect 6686 7588 6742 7644
rect 6742 7588 6746 7644
rect 6682 7584 6746 7588
rect 8374 7644 8438 7648
rect 8374 7588 8378 7644
rect 8378 7588 8434 7644
rect 8434 7588 8438 7644
rect 8374 7584 8438 7588
rect 8454 7644 8518 7648
rect 8454 7588 8458 7644
rect 8458 7588 8514 7644
rect 8514 7588 8518 7644
rect 8454 7584 8518 7588
rect 8534 7644 8598 7648
rect 8534 7588 8538 7644
rect 8538 7588 8594 7644
rect 8594 7588 8598 7644
rect 8534 7584 8598 7588
rect 8614 7644 8678 7648
rect 8614 7588 8618 7644
rect 8618 7588 8674 7644
rect 8674 7588 8678 7644
rect 8614 7584 8678 7588
rect 1918 7100 1982 7104
rect 1918 7044 1922 7100
rect 1922 7044 1978 7100
rect 1978 7044 1982 7100
rect 1918 7040 1982 7044
rect 1998 7100 2062 7104
rect 1998 7044 2002 7100
rect 2002 7044 2058 7100
rect 2058 7044 2062 7100
rect 1998 7040 2062 7044
rect 2078 7100 2142 7104
rect 2078 7044 2082 7100
rect 2082 7044 2138 7100
rect 2138 7044 2142 7100
rect 2078 7040 2142 7044
rect 2158 7100 2222 7104
rect 2158 7044 2162 7100
rect 2162 7044 2218 7100
rect 2218 7044 2222 7100
rect 2158 7040 2222 7044
rect 3850 7100 3914 7104
rect 3850 7044 3854 7100
rect 3854 7044 3910 7100
rect 3910 7044 3914 7100
rect 3850 7040 3914 7044
rect 3930 7100 3994 7104
rect 3930 7044 3934 7100
rect 3934 7044 3990 7100
rect 3990 7044 3994 7100
rect 3930 7040 3994 7044
rect 4010 7100 4074 7104
rect 4010 7044 4014 7100
rect 4014 7044 4070 7100
rect 4070 7044 4074 7100
rect 4010 7040 4074 7044
rect 4090 7100 4154 7104
rect 4090 7044 4094 7100
rect 4094 7044 4150 7100
rect 4150 7044 4154 7100
rect 4090 7040 4154 7044
rect 5782 7100 5846 7104
rect 5782 7044 5786 7100
rect 5786 7044 5842 7100
rect 5842 7044 5846 7100
rect 5782 7040 5846 7044
rect 5862 7100 5926 7104
rect 5862 7044 5866 7100
rect 5866 7044 5922 7100
rect 5922 7044 5926 7100
rect 5862 7040 5926 7044
rect 5942 7100 6006 7104
rect 5942 7044 5946 7100
rect 5946 7044 6002 7100
rect 6002 7044 6006 7100
rect 5942 7040 6006 7044
rect 6022 7100 6086 7104
rect 6022 7044 6026 7100
rect 6026 7044 6082 7100
rect 6082 7044 6086 7100
rect 6022 7040 6086 7044
rect 7714 7100 7778 7104
rect 7714 7044 7718 7100
rect 7718 7044 7774 7100
rect 7774 7044 7778 7100
rect 7714 7040 7778 7044
rect 7794 7100 7858 7104
rect 7794 7044 7798 7100
rect 7798 7044 7854 7100
rect 7854 7044 7858 7100
rect 7794 7040 7858 7044
rect 7874 7100 7938 7104
rect 7874 7044 7878 7100
rect 7878 7044 7934 7100
rect 7934 7044 7938 7100
rect 7874 7040 7938 7044
rect 7954 7100 8018 7104
rect 7954 7044 7958 7100
rect 7958 7044 8014 7100
rect 8014 7044 8018 7100
rect 7954 7040 8018 7044
rect 2578 6556 2642 6560
rect 2578 6500 2582 6556
rect 2582 6500 2638 6556
rect 2638 6500 2642 6556
rect 2578 6496 2642 6500
rect 2658 6556 2722 6560
rect 2658 6500 2662 6556
rect 2662 6500 2718 6556
rect 2718 6500 2722 6556
rect 2658 6496 2722 6500
rect 2738 6556 2802 6560
rect 2738 6500 2742 6556
rect 2742 6500 2798 6556
rect 2798 6500 2802 6556
rect 2738 6496 2802 6500
rect 2818 6556 2882 6560
rect 2818 6500 2822 6556
rect 2822 6500 2878 6556
rect 2878 6500 2882 6556
rect 2818 6496 2882 6500
rect 4510 6556 4574 6560
rect 4510 6500 4514 6556
rect 4514 6500 4570 6556
rect 4570 6500 4574 6556
rect 4510 6496 4574 6500
rect 4590 6556 4654 6560
rect 4590 6500 4594 6556
rect 4594 6500 4650 6556
rect 4650 6500 4654 6556
rect 4590 6496 4654 6500
rect 4670 6556 4734 6560
rect 4670 6500 4674 6556
rect 4674 6500 4730 6556
rect 4730 6500 4734 6556
rect 4670 6496 4734 6500
rect 4750 6556 4814 6560
rect 4750 6500 4754 6556
rect 4754 6500 4810 6556
rect 4810 6500 4814 6556
rect 4750 6496 4814 6500
rect 6442 6556 6506 6560
rect 6442 6500 6446 6556
rect 6446 6500 6502 6556
rect 6502 6500 6506 6556
rect 6442 6496 6506 6500
rect 6522 6556 6586 6560
rect 6522 6500 6526 6556
rect 6526 6500 6582 6556
rect 6582 6500 6586 6556
rect 6522 6496 6586 6500
rect 6602 6556 6666 6560
rect 6602 6500 6606 6556
rect 6606 6500 6662 6556
rect 6662 6500 6666 6556
rect 6602 6496 6666 6500
rect 6682 6556 6746 6560
rect 6682 6500 6686 6556
rect 6686 6500 6742 6556
rect 6742 6500 6746 6556
rect 6682 6496 6746 6500
rect 8374 6556 8438 6560
rect 8374 6500 8378 6556
rect 8378 6500 8434 6556
rect 8434 6500 8438 6556
rect 8374 6496 8438 6500
rect 8454 6556 8518 6560
rect 8454 6500 8458 6556
rect 8458 6500 8514 6556
rect 8514 6500 8518 6556
rect 8454 6496 8518 6500
rect 8534 6556 8598 6560
rect 8534 6500 8538 6556
rect 8538 6500 8594 6556
rect 8594 6500 8598 6556
rect 8534 6496 8598 6500
rect 8614 6556 8678 6560
rect 8614 6500 8618 6556
rect 8618 6500 8674 6556
rect 8674 6500 8678 6556
rect 8614 6496 8678 6500
rect 1918 6012 1982 6016
rect 1918 5956 1922 6012
rect 1922 5956 1978 6012
rect 1978 5956 1982 6012
rect 1918 5952 1982 5956
rect 1998 6012 2062 6016
rect 1998 5956 2002 6012
rect 2002 5956 2058 6012
rect 2058 5956 2062 6012
rect 1998 5952 2062 5956
rect 2078 6012 2142 6016
rect 2078 5956 2082 6012
rect 2082 5956 2138 6012
rect 2138 5956 2142 6012
rect 2078 5952 2142 5956
rect 2158 6012 2222 6016
rect 2158 5956 2162 6012
rect 2162 5956 2218 6012
rect 2218 5956 2222 6012
rect 2158 5952 2222 5956
rect 3850 6012 3914 6016
rect 3850 5956 3854 6012
rect 3854 5956 3910 6012
rect 3910 5956 3914 6012
rect 3850 5952 3914 5956
rect 3930 6012 3994 6016
rect 3930 5956 3934 6012
rect 3934 5956 3990 6012
rect 3990 5956 3994 6012
rect 3930 5952 3994 5956
rect 4010 6012 4074 6016
rect 4010 5956 4014 6012
rect 4014 5956 4070 6012
rect 4070 5956 4074 6012
rect 4010 5952 4074 5956
rect 4090 6012 4154 6016
rect 4090 5956 4094 6012
rect 4094 5956 4150 6012
rect 4150 5956 4154 6012
rect 4090 5952 4154 5956
rect 5782 6012 5846 6016
rect 5782 5956 5786 6012
rect 5786 5956 5842 6012
rect 5842 5956 5846 6012
rect 5782 5952 5846 5956
rect 5862 6012 5926 6016
rect 5862 5956 5866 6012
rect 5866 5956 5922 6012
rect 5922 5956 5926 6012
rect 5862 5952 5926 5956
rect 5942 6012 6006 6016
rect 5942 5956 5946 6012
rect 5946 5956 6002 6012
rect 6002 5956 6006 6012
rect 5942 5952 6006 5956
rect 6022 6012 6086 6016
rect 6022 5956 6026 6012
rect 6026 5956 6082 6012
rect 6082 5956 6086 6012
rect 6022 5952 6086 5956
rect 7714 6012 7778 6016
rect 7714 5956 7718 6012
rect 7718 5956 7774 6012
rect 7774 5956 7778 6012
rect 7714 5952 7778 5956
rect 7794 6012 7858 6016
rect 7794 5956 7798 6012
rect 7798 5956 7854 6012
rect 7854 5956 7858 6012
rect 7794 5952 7858 5956
rect 7874 6012 7938 6016
rect 7874 5956 7878 6012
rect 7878 5956 7934 6012
rect 7934 5956 7938 6012
rect 7874 5952 7938 5956
rect 7954 6012 8018 6016
rect 7954 5956 7958 6012
rect 7958 5956 8014 6012
rect 8014 5956 8018 6012
rect 7954 5952 8018 5956
rect 2578 5468 2642 5472
rect 2578 5412 2582 5468
rect 2582 5412 2638 5468
rect 2638 5412 2642 5468
rect 2578 5408 2642 5412
rect 2658 5468 2722 5472
rect 2658 5412 2662 5468
rect 2662 5412 2718 5468
rect 2718 5412 2722 5468
rect 2658 5408 2722 5412
rect 2738 5468 2802 5472
rect 2738 5412 2742 5468
rect 2742 5412 2798 5468
rect 2798 5412 2802 5468
rect 2738 5408 2802 5412
rect 2818 5468 2882 5472
rect 2818 5412 2822 5468
rect 2822 5412 2878 5468
rect 2878 5412 2882 5468
rect 2818 5408 2882 5412
rect 4510 5468 4574 5472
rect 4510 5412 4514 5468
rect 4514 5412 4570 5468
rect 4570 5412 4574 5468
rect 4510 5408 4574 5412
rect 4590 5468 4654 5472
rect 4590 5412 4594 5468
rect 4594 5412 4650 5468
rect 4650 5412 4654 5468
rect 4590 5408 4654 5412
rect 4670 5468 4734 5472
rect 4670 5412 4674 5468
rect 4674 5412 4730 5468
rect 4730 5412 4734 5468
rect 4670 5408 4734 5412
rect 4750 5468 4814 5472
rect 4750 5412 4754 5468
rect 4754 5412 4810 5468
rect 4810 5412 4814 5468
rect 4750 5408 4814 5412
rect 6442 5468 6506 5472
rect 6442 5412 6446 5468
rect 6446 5412 6502 5468
rect 6502 5412 6506 5468
rect 6442 5408 6506 5412
rect 6522 5468 6586 5472
rect 6522 5412 6526 5468
rect 6526 5412 6582 5468
rect 6582 5412 6586 5468
rect 6522 5408 6586 5412
rect 6602 5468 6666 5472
rect 6602 5412 6606 5468
rect 6606 5412 6662 5468
rect 6662 5412 6666 5468
rect 6602 5408 6666 5412
rect 6682 5468 6746 5472
rect 6682 5412 6686 5468
rect 6686 5412 6742 5468
rect 6742 5412 6746 5468
rect 6682 5408 6746 5412
rect 8374 5468 8438 5472
rect 8374 5412 8378 5468
rect 8378 5412 8434 5468
rect 8434 5412 8438 5468
rect 8374 5408 8438 5412
rect 8454 5468 8518 5472
rect 8454 5412 8458 5468
rect 8458 5412 8514 5468
rect 8514 5412 8518 5468
rect 8454 5408 8518 5412
rect 8534 5468 8598 5472
rect 8534 5412 8538 5468
rect 8538 5412 8594 5468
rect 8594 5412 8598 5468
rect 8534 5408 8598 5412
rect 8614 5468 8678 5472
rect 8614 5412 8618 5468
rect 8618 5412 8674 5468
rect 8674 5412 8678 5468
rect 8614 5408 8678 5412
rect 1918 4924 1982 4928
rect 1918 4868 1922 4924
rect 1922 4868 1978 4924
rect 1978 4868 1982 4924
rect 1918 4864 1982 4868
rect 1998 4924 2062 4928
rect 1998 4868 2002 4924
rect 2002 4868 2058 4924
rect 2058 4868 2062 4924
rect 1998 4864 2062 4868
rect 2078 4924 2142 4928
rect 2078 4868 2082 4924
rect 2082 4868 2138 4924
rect 2138 4868 2142 4924
rect 2078 4864 2142 4868
rect 2158 4924 2222 4928
rect 2158 4868 2162 4924
rect 2162 4868 2218 4924
rect 2218 4868 2222 4924
rect 2158 4864 2222 4868
rect 3850 4924 3914 4928
rect 3850 4868 3854 4924
rect 3854 4868 3910 4924
rect 3910 4868 3914 4924
rect 3850 4864 3914 4868
rect 3930 4924 3994 4928
rect 3930 4868 3934 4924
rect 3934 4868 3990 4924
rect 3990 4868 3994 4924
rect 3930 4864 3994 4868
rect 4010 4924 4074 4928
rect 4010 4868 4014 4924
rect 4014 4868 4070 4924
rect 4070 4868 4074 4924
rect 4010 4864 4074 4868
rect 4090 4924 4154 4928
rect 4090 4868 4094 4924
rect 4094 4868 4150 4924
rect 4150 4868 4154 4924
rect 4090 4864 4154 4868
rect 5782 4924 5846 4928
rect 5782 4868 5786 4924
rect 5786 4868 5842 4924
rect 5842 4868 5846 4924
rect 5782 4864 5846 4868
rect 5862 4924 5926 4928
rect 5862 4868 5866 4924
rect 5866 4868 5922 4924
rect 5922 4868 5926 4924
rect 5862 4864 5926 4868
rect 5942 4924 6006 4928
rect 5942 4868 5946 4924
rect 5946 4868 6002 4924
rect 6002 4868 6006 4924
rect 5942 4864 6006 4868
rect 6022 4924 6086 4928
rect 6022 4868 6026 4924
rect 6026 4868 6082 4924
rect 6082 4868 6086 4924
rect 6022 4864 6086 4868
rect 7714 4924 7778 4928
rect 7714 4868 7718 4924
rect 7718 4868 7774 4924
rect 7774 4868 7778 4924
rect 7714 4864 7778 4868
rect 7794 4924 7858 4928
rect 7794 4868 7798 4924
rect 7798 4868 7854 4924
rect 7854 4868 7858 4924
rect 7794 4864 7858 4868
rect 7874 4924 7938 4928
rect 7874 4868 7878 4924
rect 7878 4868 7934 4924
rect 7934 4868 7938 4924
rect 7874 4864 7938 4868
rect 7954 4924 8018 4928
rect 7954 4868 7958 4924
rect 7958 4868 8014 4924
rect 8014 4868 8018 4924
rect 7954 4864 8018 4868
rect 2578 4380 2642 4384
rect 2578 4324 2582 4380
rect 2582 4324 2638 4380
rect 2638 4324 2642 4380
rect 2578 4320 2642 4324
rect 2658 4380 2722 4384
rect 2658 4324 2662 4380
rect 2662 4324 2718 4380
rect 2718 4324 2722 4380
rect 2658 4320 2722 4324
rect 2738 4380 2802 4384
rect 2738 4324 2742 4380
rect 2742 4324 2798 4380
rect 2798 4324 2802 4380
rect 2738 4320 2802 4324
rect 2818 4380 2882 4384
rect 2818 4324 2822 4380
rect 2822 4324 2878 4380
rect 2878 4324 2882 4380
rect 2818 4320 2882 4324
rect 4510 4380 4574 4384
rect 4510 4324 4514 4380
rect 4514 4324 4570 4380
rect 4570 4324 4574 4380
rect 4510 4320 4574 4324
rect 4590 4380 4654 4384
rect 4590 4324 4594 4380
rect 4594 4324 4650 4380
rect 4650 4324 4654 4380
rect 4590 4320 4654 4324
rect 4670 4380 4734 4384
rect 4670 4324 4674 4380
rect 4674 4324 4730 4380
rect 4730 4324 4734 4380
rect 4670 4320 4734 4324
rect 4750 4380 4814 4384
rect 4750 4324 4754 4380
rect 4754 4324 4810 4380
rect 4810 4324 4814 4380
rect 4750 4320 4814 4324
rect 6442 4380 6506 4384
rect 6442 4324 6446 4380
rect 6446 4324 6502 4380
rect 6502 4324 6506 4380
rect 6442 4320 6506 4324
rect 6522 4380 6586 4384
rect 6522 4324 6526 4380
rect 6526 4324 6582 4380
rect 6582 4324 6586 4380
rect 6522 4320 6586 4324
rect 6602 4380 6666 4384
rect 6602 4324 6606 4380
rect 6606 4324 6662 4380
rect 6662 4324 6666 4380
rect 6602 4320 6666 4324
rect 6682 4380 6746 4384
rect 6682 4324 6686 4380
rect 6686 4324 6742 4380
rect 6742 4324 6746 4380
rect 6682 4320 6746 4324
rect 8374 4380 8438 4384
rect 8374 4324 8378 4380
rect 8378 4324 8434 4380
rect 8434 4324 8438 4380
rect 8374 4320 8438 4324
rect 8454 4380 8518 4384
rect 8454 4324 8458 4380
rect 8458 4324 8514 4380
rect 8514 4324 8518 4380
rect 8454 4320 8518 4324
rect 8534 4380 8598 4384
rect 8534 4324 8538 4380
rect 8538 4324 8594 4380
rect 8594 4324 8598 4380
rect 8534 4320 8598 4324
rect 8614 4380 8678 4384
rect 8614 4324 8618 4380
rect 8618 4324 8674 4380
rect 8674 4324 8678 4380
rect 8614 4320 8678 4324
rect 1918 3836 1982 3840
rect 1918 3780 1922 3836
rect 1922 3780 1978 3836
rect 1978 3780 1982 3836
rect 1918 3776 1982 3780
rect 1998 3836 2062 3840
rect 1998 3780 2002 3836
rect 2002 3780 2058 3836
rect 2058 3780 2062 3836
rect 1998 3776 2062 3780
rect 2078 3836 2142 3840
rect 2078 3780 2082 3836
rect 2082 3780 2138 3836
rect 2138 3780 2142 3836
rect 2078 3776 2142 3780
rect 2158 3836 2222 3840
rect 2158 3780 2162 3836
rect 2162 3780 2218 3836
rect 2218 3780 2222 3836
rect 2158 3776 2222 3780
rect 3850 3836 3914 3840
rect 3850 3780 3854 3836
rect 3854 3780 3910 3836
rect 3910 3780 3914 3836
rect 3850 3776 3914 3780
rect 3930 3836 3994 3840
rect 3930 3780 3934 3836
rect 3934 3780 3990 3836
rect 3990 3780 3994 3836
rect 3930 3776 3994 3780
rect 4010 3836 4074 3840
rect 4010 3780 4014 3836
rect 4014 3780 4070 3836
rect 4070 3780 4074 3836
rect 4010 3776 4074 3780
rect 4090 3836 4154 3840
rect 4090 3780 4094 3836
rect 4094 3780 4150 3836
rect 4150 3780 4154 3836
rect 4090 3776 4154 3780
rect 5782 3836 5846 3840
rect 5782 3780 5786 3836
rect 5786 3780 5842 3836
rect 5842 3780 5846 3836
rect 5782 3776 5846 3780
rect 5862 3836 5926 3840
rect 5862 3780 5866 3836
rect 5866 3780 5922 3836
rect 5922 3780 5926 3836
rect 5862 3776 5926 3780
rect 5942 3836 6006 3840
rect 5942 3780 5946 3836
rect 5946 3780 6002 3836
rect 6002 3780 6006 3836
rect 5942 3776 6006 3780
rect 6022 3836 6086 3840
rect 6022 3780 6026 3836
rect 6026 3780 6082 3836
rect 6082 3780 6086 3836
rect 6022 3776 6086 3780
rect 7714 3836 7778 3840
rect 7714 3780 7718 3836
rect 7718 3780 7774 3836
rect 7774 3780 7778 3836
rect 7714 3776 7778 3780
rect 7794 3836 7858 3840
rect 7794 3780 7798 3836
rect 7798 3780 7854 3836
rect 7854 3780 7858 3836
rect 7794 3776 7858 3780
rect 7874 3836 7938 3840
rect 7874 3780 7878 3836
rect 7878 3780 7934 3836
rect 7934 3780 7938 3836
rect 7874 3776 7938 3780
rect 7954 3836 8018 3840
rect 7954 3780 7958 3836
rect 7958 3780 8014 3836
rect 8014 3780 8018 3836
rect 7954 3776 8018 3780
rect 2578 3292 2642 3296
rect 2578 3236 2582 3292
rect 2582 3236 2638 3292
rect 2638 3236 2642 3292
rect 2578 3232 2642 3236
rect 2658 3292 2722 3296
rect 2658 3236 2662 3292
rect 2662 3236 2718 3292
rect 2718 3236 2722 3292
rect 2658 3232 2722 3236
rect 2738 3292 2802 3296
rect 2738 3236 2742 3292
rect 2742 3236 2798 3292
rect 2798 3236 2802 3292
rect 2738 3232 2802 3236
rect 2818 3292 2882 3296
rect 2818 3236 2822 3292
rect 2822 3236 2878 3292
rect 2878 3236 2882 3292
rect 2818 3232 2882 3236
rect 4510 3292 4574 3296
rect 4510 3236 4514 3292
rect 4514 3236 4570 3292
rect 4570 3236 4574 3292
rect 4510 3232 4574 3236
rect 4590 3292 4654 3296
rect 4590 3236 4594 3292
rect 4594 3236 4650 3292
rect 4650 3236 4654 3292
rect 4590 3232 4654 3236
rect 4670 3292 4734 3296
rect 4670 3236 4674 3292
rect 4674 3236 4730 3292
rect 4730 3236 4734 3292
rect 4670 3232 4734 3236
rect 4750 3292 4814 3296
rect 4750 3236 4754 3292
rect 4754 3236 4810 3292
rect 4810 3236 4814 3292
rect 4750 3232 4814 3236
rect 6442 3292 6506 3296
rect 6442 3236 6446 3292
rect 6446 3236 6502 3292
rect 6502 3236 6506 3292
rect 6442 3232 6506 3236
rect 6522 3292 6586 3296
rect 6522 3236 6526 3292
rect 6526 3236 6582 3292
rect 6582 3236 6586 3292
rect 6522 3232 6586 3236
rect 6602 3292 6666 3296
rect 6602 3236 6606 3292
rect 6606 3236 6662 3292
rect 6662 3236 6666 3292
rect 6602 3232 6666 3236
rect 6682 3292 6746 3296
rect 6682 3236 6686 3292
rect 6686 3236 6742 3292
rect 6742 3236 6746 3292
rect 6682 3232 6746 3236
rect 8374 3292 8438 3296
rect 8374 3236 8378 3292
rect 8378 3236 8434 3292
rect 8434 3236 8438 3292
rect 8374 3232 8438 3236
rect 8454 3292 8518 3296
rect 8454 3236 8458 3292
rect 8458 3236 8514 3292
rect 8514 3236 8518 3292
rect 8454 3232 8518 3236
rect 8534 3292 8598 3296
rect 8534 3236 8538 3292
rect 8538 3236 8594 3292
rect 8594 3236 8598 3292
rect 8534 3232 8598 3236
rect 8614 3292 8678 3296
rect 8614 3236 8618 3292
rect 8618 3236 8674 3292
rect 8674 3236 8678 3292
rect 8614 3232 8678 3236
rect 1918 2748 1982 2752
rect 1918 2692 1922 2748
rect 1922 2692 1978 2748
rect 1978 2692 1982 2748
rect 1918 2688 1982 2692
rect 1998 2748 2062 2752
rect 1998 2692 2002 2748
rect 2002 2692 2058 2748
rect 2058 2692 2062 2748
rect 1998 2688 2062 2692
rect 2078 2748 2142 2752
rect 2078 2692 2082 2748
rect 2082 2692 2138 2748
rect 2138 2692 2142 2748
rect 2078 2688 2142 2692
rect 2158 2748 2222 2752
rect 2158 2692 2162 2748
rect 2162 2692 2218 2748
rect 2218 2692 2222 2748
rect 2158 2688 2222 2692
rect 3850 2748 3914 2752
rect 3850 2692 3854 2748
rect 3854 2692 3910 2748
rect 3910 2692 3914 2748
rect 3850 2688 3914 2692
rect 3930 2748 3994 2752
rect 3930 2692 3934 2748
rect 3934 2692 3990 2748
rect 3990 2692 3994 2748
rect 3930 2688 3994 2692
rect 4010 2748 4074 2752
rect 4010 2692 4014 2748
rect 4014 2692 4070 2748
rect 4070 2692 4074 2748
rect 4010 2688 4074 2692
rect 4090 2748 4154 2752
rect 4090 2692 4094 2748
rect 4094 2692 4150 2748
rect 4150 2692 4154 2748
rect 4090 2688 4154 2692
rect 5782 2748 5846 2752
rect 5782 2692 5786 2748
rect 5786 2692 5842 2748
rect 5842 2692 5846 2748
rect 5782 2688 5846 2692
rect 5862 2748 5926 2752
rect 5862 2692 5866 2748
rect 5866 2692 5922 2748
rect 5922 2692 5926 2748
rect 5862 2688 5926 2692
rect 5942 2748 6006 2752
rect 5942 2692 5946 2748
rect 5946 2692 6002 2748
rect 6002 2692 6006 2748
rect 5942 2688 6006 2692
rect 6022 2748 6086 2752
rect 6022 2692 6026 2748
rect 6026 2692 6082 2748
rect 6082 2692 6086 2748
rect 6022 2688 6086 2692
rect 7714 2748 7778 2752
rect 7714 2692 7718 2748
rect 7718 2692 7774 2748
rect 7774 2692 7778 2748
rect 7714 2688 7778 2692
rect 7794 2748 7858 2752
rect 7794 2692 7798 2748
rect 7798 2692 7854 2748
rect 7854 2692 7858 2748
rect 7794 2688 7858 2692
rect 7874 2748 7938 2752
rect 7874 2692 7878 2748
rect 7878 2692 7934 2748
rect 7934 2692 7938 2748
rect 7874 2688 7938 2692
rect 7954 2748 8018 2752
rect 7954 2692 7958 2748
rect 7958 2692 8014 2748
rect 8014 2692 8018 2748
rect 7954 2688 8018 2692
rect 2578 2204 2642 2208
rect 2578 2148 2582 2204
rect 2582 2148 2638 2204
rect 2638 2148 2642 2204
rect 2578 2144 2642 2148
rect 2658 2204 2722 2208
rect 2658 2148 2662 2204
rect 2662 2148 2718 2204
rect 2718 2148 2722 2204
rect 2658 2144 2722 2148
rect 2738 2204 2802 2208
rect 2738 2148 2742 2204
rect 2742 2148 2798 2204
rect 2798 2148 2802 2204
rect 2738 2144 2802 2148
rect 2818 2204 2882 2208
rect 2818 2148 2822 2204
rect 2822 2148 2878 2204
rect 2878 2148 2882 2204
rect 2818 2144 2882 2148
rect 4510 2204 4574 2208
rect 4510 2148 4514 2204
rect 4514 2148 4570 2204
rect 4570 2148 4574 2204
rect 4510 2144 4574 2148
rect 4590 2204 4654 2208
rect 4590 2148 4594 2204
rect 4594 2148 4650 2204
rect 4650 2148 4654 2204
rect 4590 2144 4654 2148
rect 4670 2204 4734 2208
rect 4670 2148 4674 2204
rect 4674 2148 4730 2204
rect 4730 2148 4734 2204
rect 4670 2144 4734 2148
rect 4750 2204 4814 2208
rect 4750 2148 4754 2204
rect 4754 2148 4810 2204
rect 4810 2148 4814 2204
rect 4750 2144 4814 2148
rect 6442 2204 6506 2208
rect 6442 2148 6446 2204
rect 6446 2148 6502 2204
rect 6502 2148 6506 2204
rect 6442 2144 6506 2148
rect 6522 2204 6586 2208
rect 6522 2148 6526 2204
rect 6526 2148 6582 2204
rect 6582 2148 6586 2204
rect 6522 2144 6586 2148
rect 6602 2204 6666 2208
rect 6602 2148 6606 2204
rect 6606 2148 6662 2204
rect 6662 2148 6666 2204
rect 6602 2144 6666 2148
rect 6682 2204 6746 2208
rect 6682 2148 6686 2204
rect 6686 2148 6742 2204
rect 6742 2148 6746 2204
rect 6682 2144 6746 2148
rect 8374 2204 8438 2208
rect 8374 2148 8378 2204
rect 8378 2148 8434 2204
rect 8434 2148 8438 2204
rect 8374 2144 8438 2148
rect 8454 2204 8518 2208
rect 8454 2148 8458 2204
rect 8458 2148 8514 2204
rect 8514 2148 8518 2204
rect 8454 2144 8518 2148
rect 8534 2204 8598 2208
rect 8534 2148 8538 2204
rect 8538 2148 8594 2204
rect 8594 2148 8598 2204
rect 8534 2144 8598 2148
rect 8614 2204 8678 2208
rect 8614 2148 8618 2204
rect 8618 2148 8674 2204
rect 8674 2148 8678 2204
rect 8614 2144 8678 2148
<< metal4 >>
rect 2570 7710 2890 7752
rect 1910 7104 2230 7664
rect 1910 7040 1918 7104
rect 1982 7050 1998 7104
rect 2062 7050 2078 7104
rect 2142 7050 2158 7104
rect 2222 7040 2230 7104
rect 1910 6814 1952 7040
rect 2188 6814 2230 7040
rect 1910 6016 2230 6814
rect 1910 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2230 6016
rect 1910 5691 2230 5952
rect 1910 5455 1952 5691
rect 2188 5455 2230 5691
rect 1910 4928 2230 5455
rect 1910 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2230 4928
rect 1910 4332 2230 4864
rect 1910 4096 1952 4332
rect 2188 4096 2230 4332
rect 1910 3840 2230 4096
rect 1910 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2230 3840
rect 1910 2973 2230 3776
rect 1910 2752 1952 2973
rect 2188 2752 2230 2973
rect 1910 2688 1918 2752
rect 1982 2688 1998 2737
rect 2062 2688 2078 2737
rect 2142 2688 2158 2737
rect 2222 2688 2230 2752
rect 1910 2128 2230 2688
rect 2570 7648 2612 7710
rect 2848 7648 2890 7710
rect 4502 7710 4822 7752
rect 2570 7584 2578 7648
rect 2882 7584 2890 7648
rect 2570 7474 2612 7584
rect 2848 7474 2890 7584
rect 2570 6560 2890 7474
rect 2570 6496 2578 6560
rect 2642 6496 2658 6560
rect 2722 6496 2738 6560
rect 2802 6496 2818 6560
rect 2882 6496 2890 6560
rect 2570 6351 2890 6496
rect 2570 6115 2612 6351
rect 2848 6115 2890 6351
rect 2570 5472 2890 6115
rect 2570 5408 2578 5472
rect 2642 5408 2658 5472
rect 2722 5408 2738 5472
rect 2802 5408 2818 5472
rect 2882 5408 2890 5472
rect 2570 4992 2890 5408
rect 2570 4756 2612 4992
rect 2848 4756 2890 4992
rect 2570 4384 2890 4756
rect 2570 4320 2578 4384
rect 2642 4320 2658 4384
rect 2722 4320 2738 4384
rect 2802 4320 2818 4384
rect 2882 4320 2890 4384
rect 2570 3633 2890 4320
rect 2570 3397 2612 3633
rect 2848 3397 2890 3633
rect 2570 3296 2890 3397
rect 2570 3232 2578 3296
rect 2642 3232 2658 3296
rect 2722 3232 2738 3296
rect 2802 3232 2818 3296
rect 2882 3232 2890 3296
rect 2570 2208 2890 3232
rect 2570 2144 2578 2208
rect 2642 2144 2658 2208
rect 2722 2144 2738 2208
rect 2802 2144 2818 2208
rect 2882 2144 2890 2208
rect 2570 2128 2890 2144
rect 3842 7104 4162 7664
rect 3842 7040 3850 7104
rect 3914 7050 3930 7104
rect 3994 7050 4010 7104
rect 4074 7050 4090 7104
rect 4154 7040 4162 7104
rect 3842 6814 3884 7040
rect 4120 6814 4162 7040
rect 3842 6016 4162 6814
rect 3842 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4162 6016
rect 3842 5691 4162 5952
rect 3842 5455 3884 5691
rect 4120 5455 4162 5691
rect 3842 4928 4162 5455
rect 3842 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4162 4928
rect 3842 4332 4162 4864
rect 3842 4096 3884 4332
rect 4120 4096 4162 4332
rect 3842 3840 4162 4096
rect 3842 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4162 3840
rect 3842 2973 4162 3776
rect 3842 2752 3884 2973
rect 4120 2752 4162 2973
rect 3842 2688 3850 2752
rect 3914 2688 3930 2737
rect 3994 2688 4010 2737
rect 4074 2688 4090 2737
rect 4154 2688 4162 2752
rect 3842 2128 4162 2688
rect 4502 7648 4544 7710
rect 4780 7648 4822 7710
rect 6434 7710 6754 7752
rect 4502 7584 4510 7648
rect 4814 7584 4822 7648
rect 4502 7474 4544 7584
rect 4780 7474 4822 7584
rect 4502 6560 4822 7474
rect 4502 6496 4510 6560
rect 4574 6496 4590 6560
rect 4654 6496 4670 6560
rect 4734 6496 4750 6560
rect 4814 6496 4822 6560
rect 4502 6351 4822 6496
rect 4502 6115 4544 6351
rect 4780 6115 4822 6351
rect 4502 5472 4822 6115
rect 4502 5408 4510 5472
rect 4574 5408 4590 5472
rect 4654 5408 4670 5472
rect 4734 5408 4750 5472
rect 4814 5408 4822 5472
rect 4502 4992 4822 5408
rect 4502 4756 4544 4992
rect 4780 4756 4822 4992
rect 4502 4384 4822 4756
rect 4502 4320 4510 4384
rect 4574 4320 4590 4384
rect 4654 4320 4670 4384
rect 4734 4320 4750 4384
rect 4814 4320 4822 4384
rect 4502 3633 4822 4320
rect 4502 3397 4544 3633
rect 4780 3397 4822 3633
rect 4502 3296 4822 3397
rect 4502 3232 4510 3296
rect 4574 3232 4590 3296
rect 4654 3232 4670 3296
rect 4734 3232 4750 3296
rect 4814 3232 4822 3296
rect 4502 2208 4822 3232
rect 4502 2144 4510 2208
rect 4574 2144 4590 2208
rect 4654 2144 4670 2208
rect 4734 2144 4750 2208
rect 4814 2144 4822 2208
rect 4502 2128 4822 2144
rect 5774 7104 6094 7664
rect 5774 7040 5782 7104
rect 5846 7050 5862 7104
rect 5926 7050 5942 7104
rect 6006 7050 6022 7104
rect 6086 7040 6094 7104
rect 5774 6814 5816 7040
rect 6052 6814 6094 7040
rect 5774 6016 6094 6814
rect 5774 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6094 6016
rect 5774 5691 6094 5952
rect 5774 5455 5816 5691
rect 6052 5455 6094 5691
rect 5774 4928 6094 5455
rect 5774 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6094 4928
rect 5774 4332 6094 4864
rect 5774 4096 5816 4332
rect 6052 4096 6094 4332
rect 5774 3840 6094 4096
rect 5774 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6094 3840
rect 5774 2973 6094 3776
rect 5774 2752 5816 2973
rect 6052 2752 6094 2973
rect 5774 2688 5782 2752
rect 5846 2688 5862 2737
rect 5926 2688 5942 2737
rect 6006 2688 6022 2737
rect 6086 2688 6094 2752
rect 5774 2128 6094 2688
rect 6434 7648 6476 7710
rect 6712 7648 6754 7710
rect 8366 7710 8686 7752
rect 6434 7584 6442 7648
rect 6746 7584 6754 7648
rect 6434 7474 6476 7584
rect 6712 7474 6754 7584
rect 6434 6560 6754 7474
rect 6434 6496 6442 6560
rect 6506 6496 6522 6560
rect 6586 6496 6602 6560
rect 6666 6496 6682 6560
rect 6746 6496 6754 6560
rect 6434 6351 6754 6496
rect 6434 6115 6476 6351
rect 6712 6115 6754 6351
rect 6434 5472 6754 6115
rect 6434 5408 6442 5472
rect 6506 5408 6522 5472
rect 6586 5408 6602 5472
rect 6666 5408 6682 5472
rect 6746 5408 6754 5472
rect 6434 4992 6754 5408
rect 6434 4756 6476 4992
rect 6712 4756 6754 4992
rect 6434 4384 6754 4756
rect 6434 4320 6442 4384
rect 6506 4320 6522 4384
rect 6586 4320 6602 4384
rect 6666 4320 6682 4384
rect 6746 4320 6754 4384
rect 6434 3633 6754 4320
rect 6434 3397 6476 3633
rect 6712 3397 6754 3633
rect 6434 3296 6754 3397
rect 6434 3232 6442 3296
rect 6506 3232 6522 3296
rect 6586 3232 6602 3296
rect 6666 3232 6682 3296
rect 6746 3232 6754 3296
rect 6434 2208 6754 3232
rect 6434 2144 6442 2208
rect 6506 2144 6522 2208
rect 6586 2144 6602 2208
rect 6666 2144 6682 2208
rect 6746 2144 6754 2208
rect 6434 2128 6754 2144
rect 7706 7104 8026 7664
rect 7706 7040 7714 7104
rect 7778 7050 7794 7104
rect 7858 7050 7874 7104
rect 7938 7050 7954 7104
rect 8018 7040 8026 7104
rect 7706 6814 7748 7040
rect 7984 6814 8026 7040
rect 7706 6016 8026 6814
rect 7706 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8026 6016
rect 7706 5691 8026 5952
rect 7706 5455 7748 5691
rect 7984 5455 8026 5691
rect 7706 4928 8026 5455
rect 7706 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8026 4928
rect 7706 4332 8026 4864
rect 7706 4096 7748 4332
rect 7984 4096 8026 4332
rect 7706 3840 8026 4096
rect 7706 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8026 3840
rect 7706 2973 8026 3776
rect 7706 2752 7748 2973
rect 7984 2752 8026 2973
rect 7706 2688 7714 2752
rect 7778 2688 7794 2737
rect 7858 2688 7874 2737
rect 7938 2688 7954 2737
rect 8018 2688 8026 2752
rect 7706 2128 8026 2688
rect 8366 7648 8408 7710
rect 8644 7648 8686 7710
rect 8366 7584 8374 7648
rect 8678 7584 8686 7648
rect 8366 7474 8408 7584
rect 8644 7474 8686 7584
rect 8366 6560 8686 7474
rect 8366 6496 8374 6560
rect 8438 6496 8454 6560
rect 8518 6496 8534 6560
rect 8598 6496 8614 6560
rect 8678 6496 8686 6560
rect 8366 6351 8686 6496
rect 8366 6115 8408 6351
rect 8644 6115 8686 6351
rect 8366 5472 8686 6115
rect 8366 5408 8374 5472
rect 8438 5408 8454 5472
rect 8518 5408 8534 5472
rect 8598 5408 8614 5472
rect 8678 5408 8686 5472
rect 8366 4992 8686 5408
rect 8366 4756 8408 4992
rect 8644 4756 8686 4992
rect 8366 4384 8686 4756
rect 8366 4320 8374 4384
rect 8438 4320 8454 4384
rect 8518 4320 8534 4384
rect 8598 4320 8614 4384
rect 8678 4320 8686 4384
rect 8366 3633 8686 4320
rect 8366 3397 8408 3633
rect 8644 3397 8686 3633
rect 8366 3296 8686 3397
rect 8366 3232 8374 3296
rect 8438 3232 8454 3296
rect 8518 3232 8534 3296
rect 8598 3232 8614 3296
rect 8678 3232 8686 3296
rect 8366 2208 8686 3232
rect 8366 2144 8374 2208
rect 8438 2144 8454 2208
rect 8518 2144 8534 2208
rect 8598 2144 8614 2208
rect 8678 2144 8686 2208
rect 8366 2128 8686 2144
<< via4 >>
rect 1952 7040 1982 7050
rect 1982 7040 1998 7050
rect 1998 7040 2062 7050
rect 2062 7040 2078 7050
rect 2078 7040 2142 7050
rect 2142 7040 2158 7050
rect 2158 7040 2188 7050
rect 1952 6814 2188 7040
rect 1952 5455 2188 5691
rect 1952 4096 2188 4332
rect 1952 2752 2188 2973
rect 1952 2737 1982 2752
rect 1982 2737 1998 2752
rect 1998 2737 2062 2752
rect 2062 2737 2078 2752
rect 2078 2737 2142 2752
rect 2142 2737 2158 2752
rect 2158 2737 2188 2752
rect 2612 7648 2848 7710
rect 2612 7584 2642 7648
rect 2642 7584 2658 7648
rect 2658 7584 2722 7648
rect 2722 7584 2738 7648
rect 2738 7584 2802 7648
rect 2802 7584 2818 7648
rect 2818 7584 2848 7648
rect 2612 7474 2848 7584
rect 2612 6115 2848 6351
rect 2612 4756 2848 4992
rect 2612 3397 2848 3633
rect 3884 7040 3914 7050
rect 3914 7040 3930 7050
rect 3930 7040 3994 7050
rect 3994 7040 4010 7050
rect 4010 7040 4074 7050
rect 4074 7040 4090 7050
rect 4090 7040 4120 7050
rect 3884 6814 4120 7040
rect 3884 5455 4120 5691
rect 3884 4096 4120 4332
rect 3884 2752 4120 2973
rect 3884 2737 3914 2752
rect 3914 2737 3930 2752
rect 3930 2737 3994 2752
rect 3994 2737 4010 2752
rect 4010 2737 4074 2752
rect 4074 2737 4090 2752
rect 4090 2737 4120 2752
rect 4544 7648 4780 7710
rect 4544 7584 4574 7648
rect 4574 7584 4590 7648
rect 4590 7584 4654 7648
rect 4654 7584 4670 7648
rect 4670 7584 4734 7648
rect 4734 7584 4750 7648
rect 4750 7584 4780 7648
rect 4544 7474 4780 7584
rect 4544 6115 4780 6351
rect 4544 4756 4780 4992
rect 4544 3397 4780 3633
rect 5816 7040 5846 7050
rect 5846 7040 5862 7050
rect 5862 7040 5926 7050
rect 5926 7040 5942 7050
rect 5942 7040 6006 7050
rect 6006 7040 6022 7050
rect 6022 7040 6052 7050
rect 5816 6814 6052 7040
rect 5816 5455 6052 5691
rect 5816 4096 6052 4332
rect 5816 2752 6052 2973
rect 5816 2737 5846 2752
rect 5846 2737 5862 2752
rect 5862 2737 5926 2752
rect 5926 2737 5942 2752
rect 5942 2737 6006 2752
rect 6006 2737 6022 2752
rect 6022 2737 6052 2752
rect 6476 7648 6712 7710
rect 6476 7584 6506 7648
rect 6506 7584 6522 7648
rect 6522 7584 6586 7648
rect 6586 7584 6602 7648
rect 6602 7584 6666 7648
rect 6666 7584 6682 7648
rect 6682 7584 6712 7648
rect 6476 7474 6712 7584
rect 6476 6115 6712 6351
rect 6476 4756 6712 4992
rect 6476 3397 6712 3633
rect 7748 7040 7778 7050
rect 7778 7040 7794 7050
rect 7794 7040 7858 7050
rect 7858 7040 7874 7050
rect 7874 7040 7938 7050
rect 7938 7040 7954 7050
rect 7954 7040 7984 7050
rect 7748 6814 7984 7040
rect 7748 5455 7984 5691
rect 7748 4096 7984 4332
rect 7748 2752 7984 2973
rect 7748 2737 7778 2752
rect 7778 2737 7794 2752
rect 7794 2737 7858 2752
rect 7858 2737 7874 2752
rect 7874 2737 7938 2752
rect 7938 2737 7954 2752
rect 7954 2737 7984 2752
rect 8408 7648 8644 7710
rect 8408 7584 8438 7648
rect 8438 7584 8454 7648
rect 8454 7584 8518 7648
rect 8518 7584 8534 7648
rect 8534 7584 8598 7648
rect 8598 7584 8614 7648
rect 8614 7584 8644 7648
rect 8408 7474 8644 7584
rect 8408 6115 8644 6351
rect 8408 4756 8644 4992
rect 8408 3397 8644 3633
<< metal5 >>
rect 1056 7710 8880 7752
rect 1056 7474 2612 7710
rect 2848 7474 4544 7710
rect 4780 7474 6476 7710
rect 6712 7474 8408 7710
rect 8644 7474 8880 7710
rect 1056 7432 8880 7474
rect 1056 7050 8880 7092
rect 1056 6814 1952 7050
rect 2188 6814 3884 7050
rect 4120 6814 5816 7050
rect 6052 6814 7748 7050
rect 7984 6814 8880 7050
rect 1056 6772 8880 6814
rect 1056 6351 8880 6393
rect 1056 6115 2612 6351
rect 2848 6115 4544 6351
rect 4780 6115 6476 6351
rect 6712 6115 8408 6351
rect 8644 6115 8880 6351
rect 1056 6073 8880 6115
rect 1056 5691 8880 5733
rect 1056 5455 1952 5691
rect 2188 5455 3884 5691
rect 4120 5455 5816 5691
rect 6052 5455 7748 5691
rect 7984 5455 8880 5691
rect 1056 5413 8880 5455
rect 1056 4992 8880 5034
rect 1056 4756 2612 4992
rect 2848 4756 4544 4992
rect 4780 4756 6476 4992
rect 6712 4756 8408 4992
rect 8644 4756 8880 4992
rect 1056 4714 8880 4756
rect 1056 4332 8880 4374
rect 1056 4096 1952 4332
rect 2188 4096 3884 4332
rect 4120 4096 5816 4332
rect 6052 4096 7748 4332
rect 7984 4096 8880 4332
rect 1056 4054 8880 4096
rect 1056 3633 8880 3675
rect 1056 3397 2612 3633
rect 2848 3397 4544 3633
rect 4780 3397 6476 3633
rect 6712 3397 8408 3633
rect 8644 3397 8880 3633
rect 1056 3355 8880 3397
rect 1056 2973 8880 3015
rect 1056 2737 1952 2973
rect 2188 2737 3884 2973
rect 4120 2737 5816 2973
rect 6052 2737 7748 2973
rect 7984 2737 8880 2973
rect 1056 2695 8880 2737
use sky130_fd_sc_hd__inv_2  _3_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _4_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 4324 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _5_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _6_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 5428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _7_
timestamp 1698431365
transform 1 0 4416 0 -1 5440
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1698431365
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1698431365
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1698431365
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1698431365
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1698431365
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1698431365
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1698431365
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1698431365
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1698431365
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1698431365
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1698431365
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1698431365
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1698431365
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1698431365
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1698431365
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1698431365
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1698431365
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1698431365
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1698431365
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_77
timestamp 1698431365
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1698431365
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1698431365
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1698431365
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1698431365
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1698431365
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1698431365
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1698431365
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1698431365
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1698431365
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_42
timestamp 1698431365
transform 1 0 4968 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_54
timestamp 1698431365
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_66
timestamp 1698431365
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_78
timestamp 1698431365
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1698431365
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1698431365
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_30
timestamp 1698431365
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1698431365
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1698431365
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1698431365
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1698431365
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1698431365
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1698431365
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1698431365
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_42
timestamp 1698431365
transform 1 0 4968 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_54
timestamp 1698431365
transform 1 0 6072 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_66
timestamp 1698431365
transform 1 0 7176 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_74
timestamp 1698431365
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1698431365
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1698431365
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1698431365
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1698431365
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1698431365
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1698431365
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1698431365
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1698431365
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1698431365
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1698431365
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1698431365
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1698431365
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1698431365
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1698431365
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1698431365
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_77
timestamp 1698431365
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1698431365
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1698431365
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1698431365
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_29
timestamp 1698431365
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_41
timestamp 1698431365
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1698431365
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1698431365
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1698431365
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1698431365
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1698431365
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 8004 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 1698431365
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 1698431365
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 1698431365
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 1698431365
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 1698431365
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 1698431365
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 1698431365
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 1698431365
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 1698431365
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 1698431365
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1698431365
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 1698431365
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 1698431365
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 1698431365
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 1698431365
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 1698431365
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 1698431365
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 1698431365
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 1698431365
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 1698431365
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 1698431365
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal4 s 2570 2128 2890 7752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4502 2128 4822 7752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6434 2128 6754 7752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8366 2128 8686 7752 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3355 8880 3675 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4714 8880 5034 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6073 8880 6393 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7432 8880 7752 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1910 2128 2230 7664 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3842 2128 4162 7664 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5774 2128 6094 7664 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7706 2128 8026 7664 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2695 8880 3015 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4054 8880 4374 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5413 8880 5733 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6772 8880 7092 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 a
port 2 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 b
port 3 nsew signal input
flabel metal3 s 9200 4768 10000 4888 0 FreeSans 480 0 0 0 c
port 4 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 carry_in
port 5 nsew signal input
flabel metal3 s 9200 5448 10000 5568 0 FreeSans 480 0 0 0 carry_out
port 6 nsew signal tristate
rlabel metal1 4968 7616 4968 7616 0 VGND
rlabel metal1 4968 7072 4968 7072 0 VPWR
rlabel metal1 5382 5236 5382 5236 0 _0_
rlabel metal1 4784 5134 4784 5134 0 _1_
rlabel metal1 5014 5134 5014 5134 0 _2_
rlabel metal3 820 4148 820 4148 0 a
rlabel metal3 1050 5508 1050 5508 0 b
rlabel metal2 8418 4913 8418 4913 0 c
rlabel metal3 820 4828 820 4828 0 carry_in
rlabel metal1 8602 5542 8602 5542 0 carry_out
rlabel metal1 4646 4556 4646 4556 0 net1
rlabel metal1 4416 5202 4416 5202 0 net2
rlabel metal1 4416 4590 4416 4590 0 net3
rlabel metal1 5957 5066 5957 5066 0 net4
rlabel metal2 8142 5474 8142 5474 0 net5
<< properties >>
string FIXED_BBOX 0 0 10000 10000
<< end >>
