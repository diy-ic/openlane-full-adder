magic
tech sky130A
magscale 1 2
timestamp 1702732268
<< obsli1 >>
rect 1104 2159 8832 7633
<< obsm1 >>
rect 934 2128 8832 7664
<< obsm2 >>
rect 938 2139 8814 7653
<< metal3 >>
rect 0 5448 800 5568
rect 9200 5448 10000 5568
rect 0 4768 800 4888
rect 9200 4768 10000 4888
rect 0 4088 800 4208
<< obsm3 >>
rect 800 5648 9200 7649
rect 880 5368 9120 5648
rect 800 4968 9200 5368
rect 880 4688 9120 4968
rect 800 4288 9200 4688
rect 880 4008 9200 4288
rect 800 2143 9200 4008
<< metal4 >>
rect 1910 2128 2230 7664
rect 2570 2128 2890 7752
rect 3842 2128 4162 7664
rect 4502 2128 4822 7752
rect 5774 2128 6094 7664
rect 6434 2128 6754 7752
rect 7706 2128 8026 7664
rect 8366 2128 8686 7752
<< metal5 >>
rect 1056 7432 8880 7752
rect 1056 6772 8880 7092
rect 1056 6073 8880 6393
rect 1056 5413 8880 5733
rect 1056 4714 8880 5034
rect 1056 4054 8880 4374
rect 1056 3355 8880 3675
rect 1056 2695 8880 3015
<< labels >>
rlabel metal4 s 2570 2128 2890 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4502 2128 4822 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6434 2128 6754 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8366 2128 8686 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3355 8880 3675 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4714 8880 5034 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6073 8880 6393 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7432 8880 7752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1910 2128 2230 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3842 2128 4162 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5774 2128 6094 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7706 2128 8026 7664 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2695 8880 3015 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4054 8880 4374 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5413 8880 5733 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6772 8880 7092 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 4088 800 4208 6 a
port 3 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 b
port 4 nsew signal input
rlabel metal3 s 9200 4768 10000 4888 6 c
port 5 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 carry_in
port 6 nsew signal input
rlabel metal3 s 9200 5448 10000 5568 6 carry_out
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 125874
string GDS_FILE /openlane/designs/openlane-full-adder/runs/RUN_2023.12.16_13.10.33/results/signoff/full_adder.magic.gds
string GDS_START 51942
<< end >>

