* NGSPICE file created from full_adder.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

.subckt full_adder VGND VPWR a b c carry_in carry_out
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 a VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput2 b VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
Xinput3 carry_in VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_7_ net2 _1_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_6_ _0_ _1_ _2_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5_ net3 net1 VGND VGND VPWR VPWR _2_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4_ net3 net1 VGND VGND VPWR VPWR _1_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3_ net2 VGND VGND VPWR VPWR _0_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR c sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_0_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR carry_out sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

