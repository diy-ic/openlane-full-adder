VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO full_adder
  CLASS BLOCK ;
  FOREIGN full_adder ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 50.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 12.850 10.640 14.450 38.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 22.510 10.640 24.110 38.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.170 10.640 33.770 38.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.830 10.640 43.430 38.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 16.775 44.400 18.375 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 23.570 44.400 25.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.365 44.400 31.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.160 44.400 38.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.550 10.640 11.150 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.210 10.640 20.810 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.870 10.640 30.470 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.530 10.640 40.130 38.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 13.475 44.400 15.075 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.270 44.400 21.870 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.065 44.400 28.665 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.860 44.400 35.460 ;
    END
  END VPWR
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b
  PIN c
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 46.000 23.840 50.000 24.440 ;
    END
  END c
  PIN carry_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END carry_in
  PIN carry_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 46.000 27.240 50.000 27.840 ;
    END
  END carry_out
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 44.160 38.165 ;
      LAYER met1 ;
        RECT 4.670 10.640 44.160 38.320 ;
      LAYER met2 ;
        RECT 4.690 10.695 44.070 38.265 ;
      LAYER met3 ;
        RECT 4.000 28.240 46.000 38.245 ;
        RECT 4.400 26.840 45.600 28.240 ;
        RECT 4.000 24.840 46.000 26.840 ;
        RECT 4.400 23.440 45.600 24.840 ;
        RECT 4.000 21.440 46.000 23.440 ;
        RECT 4.400 20.040 46.000 21.440 ;
        RECT 4.000 10.715 46.000 20.040 ;
  END
END full_adder
END LIBRARY

